-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
l5v8Mo+oo62INcI8A4ZEAP5A8TLrIhAlzwWCdGNGj5lkcAkqc3PN/gvQijRt1259j43uBhBDzdcm
R7EmEVeHxIWP5hqinxn3mQQX8e+PeBLXz8xgIHOtvPK7N0ZyZS4jG+hVVIVkXZ5eo8h+Nv+suQnm
pQFOI2iBnHVhkXems73zahMzoQR3Pr5OFp2PD2zQW0g/+hcyZ22bA43Wd3Ggb3AwMHKWm9vOReCH
G91J5UkUOjrHTHog+hjNubp+xDcLU1Wc2uqOBJNg3Uv4Pc2Vhce2/jeTNLxNtathTvzLgC/SIwxj
fjA7CH/Y2ID0uVWXMpNXDX7eZnwBNCYxcdAwxg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
o7VghYrc4+kXj8envqWKodJ6FJ9IpsEyrltru+E0ALleYVhP+6wQ/C/kTR9xtGgC/09LaIqktMHC
q606jLp6dzGpUAErqJ5u01UaLhERVwABkVmbNJOxsWzLMiEjMO4BmIWtz3dYb9x5WLkYF8bAIr52
28TzjtWzzgFktYxgC7QDyeC2vYRWSDVNdMqUOpQ11rOI5VX4hTRdqs8IUYkKBwj9ZF0/s1lXYYJZ
9aJydv/+J7xsuq3/F45duy/HbH0B02eXMwH6gkyjq/9whBwGPswE2s4De2wMsdpKBioYUhEgTfqw
oEvDMTjiLDOWrXoN2fNMdVcx508LPEEN7DiePwaff2+Vn7jsRKHc1yPfTE84CzWBs6OFs6Plkwxl
E1OYxZH2ZcDbM6TTfwGdsXpF39Qvwo7N2T0K0UbJ0erPYFEKB7PH7Y6Rjx8pIYJXHzmnE4MQlLxF
TuXEe/q1AOUniS4EPAX2rdaR42C7y7bVu0JNgzF6bVhG1NZD9+BdE1r31/Ht5JjTU1oiLDTuzud6
mYiHNlYDolkJAgVp5QdHpQDYL+F41okt2bC4xIw8QTFCjTgvTeI8CnSx7Eoxr5C9cZMkRbZ4TlGj
yCM3m08eaYx8KAyQKO5mL9dYhQ1aQjttoynrv/zYH90SV53RDZdYmcY1EKjJNsSX5xbuFAPDfC3a
8pWDnUKVP/W2Ac2qoWGz93Z7IIn5PTjyobupqQbD2Xki1jS3+KRdV89aizPT1X6r7KfPSVQqB9SV
dmVJrLvE/WAkPMHnU63fy75Eo10kAacqZ7lOzGZnHjjGpVq/eaDZYh5QyiHFVaNRBXf+7Th1QTNy
IwdtQwo1QMh7W4G49kpLxiY34VIXe/qffMJ/O8ToTaOBUUilbxlRNyMNKIGoEOxE8WNPUvUQVP71
pW4zBnn32yZG/jyeVOpJFdHYMLq0JlA/uKPo48HhEg4qBACywEcEzBhHgUE8EP8gqv1KsA19dx56
86u8TmDCNMAG7jL9DrauFXIsMESPbKY8YQgushqxNfi/WKl0usu/YZK7OBMWxoyAGFWGGT9+/WVM
Hm9coT48+x5Rz9trfaT9PMSqfJ1q0gl0tP1WNW4ptbzgIfz/Zdb4JxS1j2zb2r1gUmwGh+IwRyKc
ouVczvhLE407uLL9CTjITZHYDseg/9VQPJPK70Prp4YFQuq/hx5d9ACdCf+oEQ9Hmpn7yiuGhVQk
bHNqvOzIxR7fX98HrdNPddallhlvb6CHXF5Ufrn0K7EPib70EH4VLy4u1lRJD3TPvgoXE4VdaIZg
OCZGlSvJa0XBQtU3yKVvfibwWgumX8CNjR+E+lpB0rvPDnOGDno8MUPiNVbmUXXb6FHbgtesTGtq
3xcwzyGWr7qjqv6KKcPpSDI7yeHxtHz3bGlxYFQzZsKV8/Xk8U3aDQSRXm3LEl/B3sXrMcAd7rHx
E8yMB3J0/bo4j5MQBt0DSj9RY8v9dXiMRAKTHeXuIaEsoawCd7lqtLyXv8QJ+QSGt4qdpCniuV8r
M60gUa+e9ewQRt1aaw+pIN0RP3Re5nLBgh2IeTC6f0fdiH6TBtAd5/r69OU3hyvhWgkxmhi2CP5A
H9yNPCno+qjjMlC+FteFPnIDyBdsyrfG3DlP+P8rLMhrcGqZGQV2xBDw/547UkSWlBFnYscVToSn
ee5IxRi120PfMSJIUksFnJ9B3lhxE1gm50/wl3SCffezQduPMfE72SrspGHxZhlSQKKHcWc3BxlH
SRa58Dr+HBNrP5FF7Gjp7KyLzuSMKUtWYMYQtBhSQiHwJc2GdrSZ5FjKtS5aELsb9E7tyH1zavH5
qyLrIFrLaMcoYKQOun7vwRrOUe+yarV4oKcYvCD9sUeBUusGLtbtyBd6EPhJroOfW9cu2UJlHE/D
COjJiEdGwyHllmaDDZsyZIDEKK0LAUrhdu21eiR4B0+TBq/ERUwc53nBsG8aDLF8AAmg6FT9pzlY
nLb0mg7dpCB1DBQ1+DJDMQx8f4s2blZ60OkzdVFTH0nmNGjozLS6K7ne9BUkhkCX6O8jfd1uRWZ5
MIzUcDoAK5y0eKDYlWoEJP5KsPtRnOrGdPXWUsJge59xKYWBTZPhmAUhlgnRzVfppUEpyHwexEAc
LCuRDkdJfjE/N+S9eIJWV3gb5DsJ3YYQGLaMGZsQO7vMnmsIdI6GQlLdOHat/wx7/s9U83U9JCtI
EGt5hYawhX1x9SZBUBp+szyxu8jFzzWvLmZhnt8aUpo/pUc1FzM3Xjse99downmWE2IAqsK+jEL9
J734kVMdPjJArA2JOjm1s2cXtNx/C6Y7ZlayY97s2RZijAcndZKLLH03YxBpGWVkt39T3VqhOpv7
NM/uLE/8DTIUh5xzeWQzfdE7ljRemK9/thfvExMGFwxynCqAw+TmnZI6fQAx1ScXy4QBlVooX6rT
GqnDJkOqFhkxQrVY5y2WYWURUGHtGUrO5HOkNLc0Jm6+yRD3AkZE6tP6Oe0oO4o4mkuSAB1OHNZU
hbAmJCJncBvyOjp9EIgHAIwq8a7SgWNHEokwvf3TfEsmbi+Fvy7rb2vFfSJHsBRGAvEu6NGjiRQP
bXIu1TL91o9i6+nMQPUygw858RRHqM1OdivGG94OzsFRfswMxHny/8CXpLNZB1J2vKR9KaBMXL/Y
ErqZNKIIvCF8UTQSAJkpfjMIMw7HKfUmobsVJDXsiQt7qe3a4mAlv18KpML155rkUPaReV/A+wh8
9HNqSOysa0cVIWBhrwHByPHxQQxB01cFnS6HjKuX/iaFRWPNkBYqvTN6ZT0unC6YGlbpiTIEj/F3
3B60zMYV3E4FJvY4tqAXRGVcamFVuINlmRxu+h0yqT5dU4BPbDmpUMK0xdzH50nYqSNC5fjZXJEF
0QqGwjDYvgftiZ8up85sy4TwsLjWsMqyA9UXaigaRaoeTLfJ91ZCUJidXjsZV6Vx3JpNkZbllr0Y
3Wgx2LJoyyVnW66+Ho1JcHh0ovbgV+MM6+XrGStjT5WGPVhT6eEMevHm42Ow5avM0YFJYUeNzuOT
M4hXyzsXWBESgDeprgaLIIzUmzEfaWrdwO4Lq3+BEIuYAqWTHfnsTdSRAZT90PcCExm+KimhMQyV
pfF17hlHev6rbTLBl1zYemSZn/raGoyQHiOFtkMDfYqV+MUAIldviVw3Sw9U/0avHVpwNVH2oQaq
1SAlspufuz7/RmeZ/drgMPOqN3xnS/GsPRHwrGfX57KyeTYINEllUl+8sKqbj6hyQfsjKrPNaRmi
7BY3IsMOSKC2xvzG79UZQDH2LSEuez5oyxbdrSzjyUwoyXtr5dAxKhwy+td6kahVEOTh2M3+pt83
/U5nwFbMBUCCcC3KMQt9Huj0a65g1eSasLNxK2wYzpusdlly4LUlxKWjgEs4I8NkWU0btOdQk/PE
i8VMR5ZSndYAqxtaGVt815Bxes/x/IOqej+Zo6yop0uGl8FwsYutj6Tw5rvXKMxlxf8HJeRASQ8o
lNgr64JXpIsNqqZDmbIAWJhjCp8iNXIGrul20jit+dTXtnajK8AVpyuPI5z3OcK6lqibOrHSiJyZ
pUlZyZR7RMyQOpezvyQ1MKZcdRStpPEDi80zEFQwP1fkPWtBsJQoNmdQ8whxGCUYCU9ta9yyJxb9
rMeN/0xpmLhhz9iPSaGbV0FHnZsw2y3fCVv110DMpfcdnEVarYJQhEjP2wPN2xIC5oVqD+oiqnqc
neeF9Q1SsvqVtDrm7tAAibHNkfvJ9SdPF4JFcdbOAqxG5eDtrzF3e5EdsC8A30fJllzSO8Crhg1O
LD5/ZRhaqsZFrb4EGZcRUqoJXYrdGcmx70B/ShtFZIfiA1Vcz2I5TXaEcF0N3nuA6thOiNv7PCHv
0XS5oVc3pCL85k2QD9U7qQSB0IKVDJkgTeBhoHzBYSrb2sbPkXNGlZOVRZftnb5qJLKlLRUlZwoP
DleI1Yxnk5UBFOwBZa6cg2gLposXG6/EQeLPN81Fipd/jaj7Nv2lVPtxbT+NOU065M0Vppv2D9kY
pLMo4JaY039hL30QPm4Nl/f5nViSE2g0U5sJBaB3ZBDA81qHDk1Rz+Cw4QElsMxHjbx+oRY2gICI
KiXaSkVhYBA03GsL2C4ZffzOkcGM/+LguGsGo3fgMgGRw/moFy5r6M2tYxOwC5hV6iSdH/T9H9Y2
R4Ia3HbYlTMM2yx/CHOf/OsTU5AXwBdXIllk5+WTQL4MNDLXFe3rs3PzZ++Sv+T2EBmslycoyHmh
Q6tQI83Cd6PkaRnjpjzMzII4uw6qCX1pq7iJUFcahZMgS2hS2FhaeVITlaTEKGMvTRoGEW5DXGEf
Fd7SG5GfjrM4bxJSOuKNNlPXpKFgV+y3x6zkr33Ine+g2lM4amUtvp0xdaGhxT5Pi83v1CBbhIwl
5vb5qb7ekupXUTKqQ++fzMXKXV2t3M23diMcHKt1g+Bz4vu3dLUQqTKGC8lfZi6uerxttjkF6jjj
1Hx1MFUvA6Wc2QcYw7bk9+whw2q5BCwv849EmjXEaw6N/uXHQHOyglYObQSykQ/+7kufOZZlL8ma
ZIVnqUGVczlMUUDBgdtVQfb+NWOL9Kb2Ao9YuSX9ZnXFnU/L6crhW/fy0kJiLo0p3GhzpaTfIHn8
QsQadFl0h/2J8wHUW1YklcrOb7FanMEFPazEQWPTzZNJLK6Y+6V0t3S3kBfp+jUwPZoNshOqC/Vx
khR9c1FgBm0uNLlgkufukgBmfvDvdKvGxA8F/NXl6U5akt4dzmW3c6t5vuSyR5EAzi0Wg0mzpPSo
jPxtdPGF+oLSgS8uUsEo9AVJIvtn2+jRIIUy2T0ccCVPcioD/3n3l1WDCdgm79tfENTNe0FMMnzc
EQ9teN5hSHXlljh8OXyH811eaJtzdOhU03yeAW0TORC5Ms1658C8cieBwDZBEyIZleR/MBzGUXim
+g4tlfj6bHj9OfY/U+Nt3DrrxQFLXm97ZAHrIhIi3Ip5F7Fz66ln4l7acrsuRAPFfBdH0mDiib4m
WBmEXeumyJscti8FZKafuvkNigHiZr0qDJ1RxMosjBIn6sWsFerBzl/ZFhaj/THSbJchulhpFoKz
jF+QXz4g0hcaQatZbHms2pJeCi5kgMN6Op2v6DehYtJcVKgvBIYfkNol37Mypet1E1wt4YC66ZU4
zkz7rdXUZRvFXk8Pad3JFEqKsn+yDlD51LAU7NwTidC+CL9s3o/+vXER1k0hy0V42FhEII2BcmzB
JrhYaQjmsHTpiEjKz823Zq7S7oQ6ZVpZgFh4uLM8JVZaOAfreCusgU2QaDbF4pn65DfJf4fc89Hx
9txFxh6BMS3dEh/mT8QPI5MGi7bxrcN0XNjddxg2OjrsGzgdJu5CbvIRxOaI0/LfmKihRhxSdjqd
FSLjMK6FNAZQs6Ak9l6wqmnxr2hADqJ5juOTSzXlM99Inn3zt2Q2a9RyNohQkzStoIixF9fGuufo
y1euE61sRJFtb1jy8kBoBbcrM2Vc5oO9aU+JCNmThM9+QaFrX9Qnvnw3HQrLONc5cNFxbycsb1DW
c1ZtKNKhDQ256deVgARUFqaWQ4GojLOLO38uNQkHY3mN/GAHeX93KdbKKMOFn+wybuMKse+F2NPn
gEI+nKyS8wdRe2e+wnwJy0pG4mVxfgu52LShs7w0eX5vzhPL4nuLn7xmuIbPBiRWiOsvSpnM1+kI
Wf7Ixmtgjp+6IE8TDMBKGgYIR9osfVbyrpjC5o94gYqTBdskpPocwLJym6TtF5WDfb4F1+hSoY4N
F2/bjtrDu5DH2uKx+p92kSdvtKL1dJ/Ip2HHax3CWAmDA+ERimyxI0rZ4cuqfvOK01KUeMwcUlm2
xCHFy7VkHo6l/4yK3gd9gjj/HEecJwLiXxQg2T646h+XzsUGEejzjIzLO9+X2wc+KKf5FKiyqvy0
nud66QccePXwT5kgbWYTcOzosJidQZWH1v51RzMDTw48qHogjdaxU4fQbudGYrZ0Ng48GLYiaau4
sLUHCu5YiTaSZmEJ/KKuh162IrgeF111ZilWWjnicNUcRgECyFZbAJbQTzHEbW7/wheRBR1jX0tc
F0fcZEUr3I/MaW2Ad17GOPbrGNb42VFj8mxPGPmiACbsDMMbM2JxD5NHajnm2yKVoVN6NrAGSueh
qfA8Y6d2Vg1mrzZ1aYhc2GwrvCwaGStUUeVR4TJu3+nofCHQlrxU4Pt+YnELpNuplARDBxywIZ6b
3FmDWVOtSEx3/3svWER9lXl8AQjOLsR8qVhnAGFlHUER3iSoX9YHIfYrr5Z4DUJ1xeNDWFUKYXD0
81Kbhp0x1xT6yt0+Fi82ffQOoggJIzO3v9WowPyKKvH6HPbi812dPnjM1RxQ/H0v0xgqJyDMN/hm
o4N/OR9aTDZSbuEo6ubAb8OWzmJKuFoI8w37s/tO+bRI62lKDH2CMQos1uS5wrCM+44SucK3UZar
h8v3nHRNXau6675d2Mey7pL5VHKq4aWqHhwEt2e4Jo1jxjkU784Bv15dr9snzjnIlvQHECvLn2zh
7xJNEc0SQau1MyzGzwzrS26UsAYERFBKHd3hkkLidxmURDQV9JLQReN5DKnf5DiPYzNiC0LusIMQ
D9dO3SNQpCgZZsXrC8xiE+B4H5kbYHgESc7eDwQwQgKxmygM8Q+5zNWaLU9+ieNlJ6N/+s6fA0ew
UVMb6NMsxZULHqCMX6beqI44akrxt48nq1hfsiDj5YuU52KxXELSKXUdKUhIv7NkuEG4MI9nj/fc
DeKiueSqSb0702xhL1m3BIBsZW+FPQskCQ8xMOjJULCYIY/KBtqeqFPoPdljk7YhD+/ARlrrag+m
peXAK6ORYN5BbbEbVxDptdX65YuYRoYmL5S1qOHLrkx3jn/9sAeLjN3yzcxXNtX3WUCQ9laRZPWu
jaYLQvSkfSfbXYJxPf7KxWjKV9jVF1jgRozgKXde5DbQwcDM417PX8ckPGBmJf3/3Uo4zgfNiAyw
6Yjk/2aCFFurm7Lon6e+Wv8WYDfd0f77Epe8vLee+f/gu5AU6O4aSQmgdh5ESmF1UHIpiA2oSdvQ
+m9QAE/+Tyi4QyTDeymBAnR5iWfEzDX6gs4V1ESu5xgvhPTsDPw7atDi55vntIkhibPbWk0ttWha
ir4CSjINA92ymhtJK+o2IjadBVGjdNE2T7cv2V8HxftO/9uMmOxGrwenM0Nka4b1pA3ZDEr95g7x
OBMtMcMCQrufZ1f5T4pj/7Em3N7HKspUM7MPjW26tW3iM0aIyodc315DGp10+H4M2xUXO1UZ9E0N
dWU0lhGz2Zs2rLbVEKOLFDZGQwTPLdqUDA3YKOsId0j5cU7X8mGu7RBiNHHLTQoBArWFjQIe2POh
ZFnf9hTMjkmNNmbTDA35oFqEDY4ynY6QNR+Fz2vSLbl26f72dcbejPmrbB1I7CIfkZyyEuGMOtP/
4rRmFznS703DwmspD46qAVO5JIDS+STGrP0c//STmR7rkgGTdpLIE6LOaTlSLu5whGwTp6LUBJCE
ocJajHMhxP6h1OShgTNeReMsNNl+5HkBCrMYbhVxBhVGtBzwPeagprhgpLX/dIrw4gx9PRyQPuPV
9GeZLuuzqU/U0xxnxBE5tMKZtAFRqp5FNJ3Y2XRfV5d/N1BVMi6e1KiHuixoPMZm+duYr2FuP9ur
G/jQw32tgbtBdYXkLcj5xkzt2EvGFwM1MHHaOpm/kDhCfLMAcdjhLKoOu7bW/RpX5vjaxYuciiUp
FhM0jVXB7IAp4JlF33fR8c8D0CZeNwg+q+UOuSMWIJ1uCLIhySqwugV1ULRlEknuuOPR8/O0JlOR
dU6SGLVYnsk4feRzX1dWerFz+smstBlKwLvHFUXVj6olIJEVbiYbHHYiZnxvlv2ZopUxJPCpmqEA
MQ/zZl9kmeL/lzGS8OEkyDfd9D/iK3OfaRhLrV3LKvxhKRC/I3qNLDv9WWvD26lg05P7SY62sNrT
ZcL2u2uaCc9ASTfq7tAWkX0gW0o4F6S1yzYGSn8DAX8FJeWHbKNIOp9JyiDE0dg3pNTYuI5NT9YV
NvwmhHl1w0su8Sf7UnaoPVOlS57cVEwkmVGr346vpuEMQIEH9ZQTKtItRpkTTQ8W6ZPgwelXof27
6zdU7odmgRWDgDTathgsdFPUwoK2EP82e8Q9eIiSGPRUr4DAGqZ8hmDKeuGqmu3ROhEDFJ6JXgvB
5oyfchlas1SGndoJ9meY4esznrC8LwOmBixDen10vwc94KEuq09iArlqp9SvsGOFE4E6pF3tps2Z
o4gBS3N+4RKm5b/0IxqU7mO33KhuCNLmK1auPCAMiKBraLufpAORfb6Htsbaf4siCAY8gE31sLQW
5yvwMdF72VKz0x6S7Sk5lfumTTdQwUiJpppDCjNjJcVQJz+rdShwvF3Owqulwwuu09J4rOfNtb5h
2FnDO2YezyNl0/UNqUYqnFtODFHoerCfLDYhZ7uEWFNtbnOxDho+7TJFoWg83u6PjRVGQzWOpSLx
oZW21n6U5/Kwf2ANeizx20U8gzt/w9sCvjaE7Z6CnneFjEcoHdZysoX7g/4GjKH35HaO9YlGcrMZ
pxlFEZEJA3jsuj5gYmq2+kZL9sMnqCEnwpiw1vjjEqPTMo94EK2cw+FCNTKzY/+KDcA2xjzvyGH7
GXoisDVn7iaU4qVpPziw/gfyn4HDooJvlzbofbD8cEQLksPxTPvOE92xx8zxVsYqIepmvaUvHXSk
gOeUtEgKw+nhLR9nWXLbpdtQ6LFKLObP8uaDVmAZG2up+3VAulIWdMHbxSze9P7gZBI94TRacKF9
VCCnThpCYG1Z48EslryJkhnmNWY/XFd4wDiQ/k4pL0+tg24YyL+9AmrMK0+IlSxOx9/nHr+vrGzm
vGJWfHa7bpcIe/nJOX5hEn8KH32ebMgETszcuWsZEI3HQZYlTLhZX7veZBMGCl1pQNFVqwDCED1o
lKoGDh9T8zvD6FXyr+9/eG0n2FUSUx99FKfVAzbWPFvbTUoK9R7ahNjO63wEe/jgjpGSs+r5xxbF
Hnaoz9iKfrmsjLc/rhAINtGeAaCJT9F1cPBaI9PVuHDm8IcNZ97HZnHicLbBCuMni2amDlW6LOZI
a0c6SrA8UVAt+Rc8S9CcN1c6wPXxdkgimHLV8n5h4xaJzwhUNEpGHOkVi+raBFt8jJ8LlAtFcf/5
NjFLAKTkbl0qEOvbaNsjdN1y5nIKPRqOwZWT1HvRNQ7MukwnAmJcikDPVcyrqGWE1nFbMVYfXIB/
2Vd5wnXqy2vKGigtKElIAAF7UJYhaS4sgcK2b09Ql0pjr6mfnroOeqRCwy2mcZAdzGOhMH50y55g
QzjbjTwzdiVHEF0GETudVSv4Zs2WKEMqIl3D7q/KnnoWYt4Ti42IgQ8Wkb0oUWUKKqYywbPfZ2nq
JxYdcos7VhWhzllWtnj/kKEA+aENo/DUnq61FV1M19I58dYNsfEFM0tjcOboHYS3tmlpfmRVG1U6
BT606sOCO6jHdpwJ0dCM+OmEbYBIgKky5Xz5SaTmPLWdT1pcBvMp6YVl7rBLKTRwynWRsQdAQ1AQ
yC+ga1EpRAyEBPD82oxg8roHJK1HNKGUOcKSi1s9UXIJJRkHGywfCxXJ7qvuRaTFXd8v3QigsSzl
3MjsTDxmSj6min3XWX9DjHs0PPQrCLWBv9Xm/lRDAlYnyNoh1x/GhJrZP1RrpP4o54eVsOW9EOD0
f28iiZ+1BDeZmFKYD+1maoSbOr2VRnTUpvCLlRfxISD2KEC+iRqGtldylKUJtOH+mGFkNN0dkVZA
OK/o6rMiwFPhO7FgfAOvHeQSzZXxIJq3BGE1duXHGObMJytrNkwml5n8r/XK+Gis3OM9L8hIGV//
n17BZwp2DePR8zhdAgYjcJOFbAW1qXH7Ceejla3L6+c/EhqmWJqjzkkxYWVcvSAW/F6pQc3SmN/n
hcG+yRO5zISSRwwerH/QN2Cy/j9SkIQ1GPEBKL1SC0Hy86BHQVANCaRMoAtBio6gbduqXA7/QUaW
ZkXg07CGHSbOrfSU9FAemDEAQ6euryaFRtyDLVEGVO1WmF1Z7rya5XVJX5mOLeMhOTV3coxkPwkA
THBc59peBtwW5bHBTHPdjP+b4nWAuozSfYpjHKM6evnoNk/xb+nnXlqGSw6hF3ce2VdpJZjq/T4r
zTNyA1Kvtvl7XUN723y38R0PprzCr1/AqjLpBs1swrmGTGn/bIZKvoITmfjhhdng93hxpFe6ZcHm
pdBrNE/dj/PCPy3c8lXFgkx9IINqt4/3cgUU1mTeimj+sUtLLl+uGJ+3CPW8D+C7iWG4WNme+ViB
FfSJrEwXpidgKksxPYSsFokmBzoICnyrBeretly2lLcvB3HPD173maVYTmhoSxX4JSSyUzgmwzI1
uwSFQI6v8NOH4IlLqYWq4O2DPKe9lYb009hLQ5Mq53fBP3FrPt8y7Llj47y1dSMsjorEY4sConSK
b+ynF1FQO0//RjgxWMv/6QryBE70tUyFqfTesxoq6vnWuOEc4IZq4Iit/A+rJ8D6G5u1u551U+A/
eYKn3g2gi/dcyVq2gw==
`protect end_protected
