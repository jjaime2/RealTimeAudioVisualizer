��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S����%J�b����j`)�u�B2z�l� ���#�p7L�7>J�ו4Ű~;�W�I�]�Ec|f�)s��˓ߑY�u�����|��
)��0fkh˔#�v��b�ɸ�* ���g'�����3�93�w'�%>~07�I�%�E�v�+J���q�[���s"k,B�ɀ(L`C��E��"�*KEBA��y��g���$�~mFy��X���x�,ᾷ71mѡ� �<:% ,I��nu�t`���Om-хb�:ǬۺJ�:��\j8\�(�_�Fq�֫8�+1o��3�p��]��ۄ�Ұ�"e�0����G
lX�y������ͷ�TQ�' z����y��rG�b�Wy����N�
b��W-ro��7yΓݬLw"����T#��jGG��BJ��d�]$M��*��^��٤�c7Y����s.�ʍjf=	�pE2�e:E%d'j�Aʃ�,Ą����C��a��V'�;/���������M�����K,��?>P{�\m�㰋�����PX���e}0r��`\�簸�S'��*#�d����-�׼/� ���KP\�#[��"P@��$,j-Lg��� ��$"����T҆2����s<����n[��&����#r&�/d.���j�!7̀�\�����}7"������z2Qx��Ya�a��_��mT��Xe�H��r��g��y8��p�&���GY�A�hA-L�6��Hԟ���E/�
k];�0d���{n�P����>���iQ]?�R���|BGdڹ������u�����(�cGr@�lݽ��5�^�*ѹ���M[��\�!A��gs�#�W��sݳ`oxN�6
ق�6���m��nMo���-Y��0�+gM���n����8�/o�1�����l,np>��4��Cc
Hj4�3~dƞk>����^�������磮t[��)�n{�Co�?c�ǭ���޷E	�7G�F��i�!h ��&��S��68�H�p0탛u��/��ɢK}$�B&�qڸ�H�]�#�O�"
)��+�hcocC�<��J��,��q[�FZ� ���g~ˢ<�.ۻmБ�1s�����܌
0�u��"" �N�?�Jɛ�n���mբ�T9�n�·hld7� =9�C�C<�A�#�'b����zT�G�"Q�pY�t*p��Y^��S�@!Ue�6Ts�هcϐ���r�ъ-�~����o���<�hìci��	��tGۣ��a%bٓ���|�za�i�E�F��xt�9B�u�����T�W�6=�6���n^��*8��f�2geġ�=w�V�b��s��� �%y�x�
����6�#��:��/��H ���>W�������w	�Ԗq7hdS�P��D2-PZ������H����pS�Y� �z@}������:�TS��S{�1ȗ
yS>��D�����p�Q��)G���j��.����;g�a/I��Z�{tA7�����[^dm�=aط����P����7V��N�!���^J=��׭Q/кIQ^��Ckx� d���(������rW�KP�3��J�����!�!s�O�O=���DN͸�\�����:O8Ѯ���^E����'��-�Oh�>1�G�0uA��>d@�7�?:C|�M\��ڤ <:d�B�+��@��$�TF�ҵ	B �P6F!�&#�,��=t�ܧs�}��\�(0q(������bn�_>|
���f�n�;��)uWXΊ'�Y���LBJ����꺽^2J��?�R^�����G-Ez����6�!�|��G0���Z7S�?�P��A��fRsԘ�0V�ZX���,��\4wl��4{Ͱ��wв���1 �#o�;����u���������D�D��bqۈ;+7ix�V<��XRA}�C�����S}6���#�|&�h�J����>B�2��R��=Ȗ�8�k�邲��'	��b��������B�Fws򆱄i�]���y��pš�d�U�|��ho��R=ӻ��8<D�P��vȇy��Ctv�'|�}�Y�kE�5�t�^b~6�\ ~J_�h{��bl�;�]�B̼�n�^'��Ҿ�=�r���v�!�a�;=�3�?;�9È�8V���.g��%�k�E���eBo9#F�q�]+��<":�x�@����[t����XVh����%O����T����چ�w�\����]V�R���]���0YǦUx)n1�F��E�Ϩ����ƹQ#��5��	�
�%d��yJ}��������M�psh���+>�@#o$�	�����ʠ�'Eu/�	Q>���ޔE�k�Kk����f��G?�<�u⡺RJ]�@�O�P��&�͋��;*�]Xƌ�^q����	�O�P��>&�;����9�t��~K!��L46��^����\9�����D�%�����e݂�\=�?R����53(?Uk��ME�Vi��}C=�`sVw!�u��(l;���<�0ԅ7��������{�S�pW� �B "f׳09s�Ȩ�x�{B5?�#VE��o��T��^x>�qN?������͕�)
m@�ғߗ(��JZ�&�,~2k6�_��>���_��f�i��aH����Yޢ���7���gp�n4�yZ�?�ǆ$P��dkz��O)�+�:�Nj$���r�7�G����,�m�V�&�mMӸ	L�M�lA��l�D�{���l���X��I��dG"�wG��cObșF����Eװ�Rն��ݱ!�`��e+>7΢=�g��A&C�6�_iE��a�d:�ru�;��K�ՃN�)qlm2�=�.�����.��ԙǢ8�	��A�>]���|�ܰ�15���[Đ����C�r>%LL=�/ndSNCh����!��WW=bO �S�i9U, ���@�k&ЀF���rZ�������sdi�Iу�YH�Û'BY��A����j^w]�J��8�I�,/90����h>��L�!I읔������X_O_������9��{��=�'�V�S�Yv�r�=*G�V/�-x	��k7�%4#��Dc������W�Ҵ��wN��vж��Қ��,9%��0�#�U�c�\j_��+؉�B�y�ݠ&]�!mh
�7ծ�e0H��!�\t�?W/����JJ27�o$�ԁc���uT���U���~&⩜�.�naq�Z����U����<S_���4"m�泴�C��Ji�K.L�}=���3��((jM�yyw��0껈ԥ��E��ҮF�A���X���)�B�hɻT$�x�a\�sg���R���_��������c"z��P�?̏2�fz`��s��W=B�""��H��Y�.�����>�kK\:��C ���/I[�(��s��YX�l�oh�y���5@��lu3�� ��U���'Q����̃}\���t5!�ORm��9�	Z�:�xH��Tl����v.+~T9�C��(S`���W@��]ԁ�7i�W���/��·��3h���od2�즸�� ua1v���%���*jX6c<=l����:�	GN�2��\���f��%ʲ���}�9�`�ba�+*����]j^;n(�Fܞ��W��9���c*.cfJ�V�>����Ea�Hz�eNK�C`ҝS�]�c.�\���
�f8�gmƛ7�[���[8oL���^*�.� �6���P��H��OP�C�#��2�A| *���f@	[��O� NSS탔0:�z>Fk��F\)��d�H�z�pN�ǁk�EUf��E��OW�+�Ty��(��\�`�B��TV��8�?�Mq�s�L�Ha0 �mlu���'��J��g��hy��FCI�q�r�u�c�U1w0a�a,*�+NH�h�1+?J�|�)ɕ����L�Q+�Z���h��aB��-�d���cԌ.QBR��B�t���?(�5��T�&Ch.>��}b�Ңg臀y���M�r�cCXl�Gk�q���r4���`�L��������z_L��\��<�HX��ݍ�z�b�W	����jd���w�`���]KU��D)Il���Ѐ�\�;j�*XI������V�;S��4���7l],�~M��T��S�-D�kB�_qy�⫃�h���I�<�5�Ve��Ӧ|N���n�|��S丳3�;4�=��_fwn�ȉ�t��>�7YE,�� ��A��#$y���L���5���(��}�҄m�/]]���R�($��0mɫ��zkw2'��Ὓ�q�p,cg�x�ّ-�h�s ���� -��Om��œ�B�1r���+�Q�A��Ԁ2<&
�r��"�Z�s�{a��ut�����Kjg��F���,��R.V�^3l�0i��K������`P��RMB�ذG�M���"������z����RSe���*���w�-�;z��-�-��p����J�!g.�K�J^/MnW��p�3�6h
��2k(��d�h��v� m$n���X_��]CwW��ÿ�}w�0��-��X�:+;����$�|K�*"Jt誤"Y_ov�蓛o��Ci�����q&H���]�;z�	
'������L�%_�G.dŇ#I��F�^#�XW+u� ���Eh���6B�:���.@�;&�U�����'�/�gr�^���'m��I��xQ��1�kh��2�b��ԍ�?K!�PG�I�ۖ��hjA�.���R�	���ǐ V.ܩ���P��eV.Dorti==L��	(��@������L�Y4Q
z�#̣�X9o�Ԏ��q��&��V����W�
r�U	�h��+aK0��=ݞ�*�������&��>�u,8�MsA�)�0]h�����0��Zܢ��oy��~ ��7�ewGE�p�\����NĿ3�����8ItT0���L�!��+K#_T����8wE.�K�� �h�t!��/p{����	-�jG`�.>�c��I;�s���ៃv����KnGb9�C��Ƃ��X��6�YU%Ar�9Ҭ::�ϫ���PJ������K�=�Xt���¡�+�GF����f�E�yg(ڠ�J����e�R%[v������B�E������y�itb�� W��J��Ώ��'����$�"̱dV��f������o�n�fX�vҴq���X����~1O�ϫgm_���6�X��_�+�Qjp?IL���٫�UCr�!o�hD�}���>�7P��[Zm#�ݳ@���זp���o�_QIC|m˜A~d[��+%�uwܶ�J܄�7�TA	�49"� 3�uZ�}[ ���3-�g����2DleI�	М7�NȎ�VX����*���p����� ?�
�V+]�bl�\Oi"������C�ອ����chn��e�����٫i�b"K0����N��(OG�'����]m����Qu{���F꧘6����P�����y�Rl�*�oH�aNo�m>��^ϕ!���KaNX�wE����Ns$f�_�,�/�l��}�
xY�a��6�$��/�J�U�rlq����u�TKZ����w�CO$�q���B����%Fn�=�-ZW�v�߻%MNC< �el����kk�ܾX����l��豕�-��s���DD1u���O��3���~Bl��2�\�QC��_P�a_(���y������?
9�t��΀�m�u��r��g2'љ(�=>u��,��Yu�X�?��c�SԢW���1�:��T ����\I��*�� �e��0p=�X�2E��#^�ʊ|X�pd� 9+�)g�Q�E����Q��F�vL����a�l�i��G=[��F�|y��&��_����{t�i�T<�fY�&��g�"�	��!�P���J���}�ƴ�zŮ8}o dn��7��E�N��(��b��r��4	ZPyꜤi(�R��U�P6�tC��AR7�{ҔK�B�$k�l3�<q��N�Pi��6�_��8+ڡj��O��YM

��	�̠�|�]�3�����n�ʹ39�ˢ�'.DX��	�榀��6*��`	��h�!��H���u"��!���K�	�Щ�O)���,���╚3���0�uҫ��[۫0}�?�v�"%���0�o��%6��4��G��O��Ry���Ʀ,&�
ȡ?���n���AQ���s��C�ygz0����;É�����ΑI'�)<.��8_@�UҶ�J<�n.�I�d��~��.����C�Ը^xR��R'���ۉU�D�q��y�'�}��);��L����D�ľ�zx���W�J�Y�+8�|��2w-�k(�/;j��A�-WOt��_�Y%�@P-��T4t�p)�b�����'�@/p�Xk̬�J�5)��kp\�Vw�������6��;zn�ؙV ϻ#}3�_���O�E�n|t�|�oЙ����D)H��jޯ����3e@l�p��!��o�Q�蒹���B1TRE�z���x}8{�c�w����?�N��Y3`�� �{4j��Aj?���U��{��F�[����3��E�J��8�1C"T�x_�v7rui���m�ۭ��
ۓ�硎����P:��E�]��x��R�1���l�����O���
�һ���e�F�P���u0�:�A�D�q!�+�Њ��ޜa����"�G���_js��q�%I����$� N5vc��ؓ��W@�^T
��Ͱ��Y�C���%KCF"�6s�aְ �d`U^F�f�Я�[X��dG��}����;�mn�(��}΢v Z�e��[3S��slnJg�(:M�KQ�bJ���]{�k"Qo��-�T���ُ`��Zs�=O!H�2i�pnDn�c��j��̓�-ep� _@���R�Ϻd��;�m�(��� H]�9OSw;a��l}6�!ց������i�m�t�����X-����=lxر��q�����]�r���3`׸�Q����\U��
a����P��GVZ�,@,�!���<����rw��AFu�!�(]d,j��؍�`_�gZ�^��+��R�ܾG�Ni9�����YHG�-��G�>��:[�G�7C2�6�n,|�s�q�J^���;E�o���2�;_	?)���ѶJ��E��}�	�A}��śk��+"l��T�ٿ�>�.q.��+=B"�zx+�0���ؒV�޺��w�w��7��W(�t4�?��0�:�E�e��sex ����;�y:�Gfe�dt��I>�FJ�MX��C���0(��篨x�>��Os;�~��,�
������;9"!8��Ď�����m5��Zk\&���E98⊋+x�	jf��^, ��ڤt��@���������n�dw�� s�ZJ�nBZ���(�8�M�U�=My�$�[��i0vDo>�*֖$����',����M)wŞ�&��Yt�8�.����.Z��"5�e�.9���hO�!��>u����\��;4�{ٌ����R�ٝ{���iPN3�Rб|��o��X�`\`���R='�=A��@i-��`��J�B�3��S��Ym��)Z��z��k�Z�t��j�K5�p#��u߾�)��\�s���׀��_;V�%fWz����K��#��l�.A���|��`���0��J�X��߼Z����њ=��37�\+���N�K.�X�C�*�`s�M����r�!R�j-{����dV�U���̾���o=hG��4��^�}S�.��Uf�z�7+˯N�0��n~Pgz@��yI�c��'�6+Q�|MW���B�-���Ί��5���*=�qIKL�+��ٛ`���Ɍ}�vf-dX��~��<=x�;~ݡ0�.���//�/yx��o�v^y�� !�I%�-b�����TbB(��ө�J���w!��;���PQϷ�%F���:B�c6�q�
�R[9t�F�� �o4ؚ��c�JpA1�FlPMg�n��r�,y�ȧ�� i�%���$Qd�� <�����쏏��24Mϝ+�L]~�
���?B)������E��"Ư�7p��(������:���$'��!F�w�x�.�s�c���5W��#+7D%�2�$�?�ʻ����� m��!�*ϵF��F�z��z�T��1{bˏ��>$�p��[���(��n{R�O9���n��+���O��F�� �;� �4ru Υ�iX�qZ�{�Ŕa���F �l �b>������� ���l_�i@�C�Z�v�+ �8J�y*�]I����%�8�4i���j�{�v�>�a8yy�ק6������C��r��}4�mf_z��^���C�f�ᇴõ�K�[~�õr��A���Dg���@g�r�Т�uP��,8�=���h����@|�"��~�)�Du�bWsP��Q���`Nx�8�>�nU�����!�3M	�G���<~_ݿ]�m.$���&)�
�:�3��ٶ��+�9����)gq07��DM���O5
��� �2˸��@�;pld@�(/��Lf���p�)����g���]�"��'�j2g L94ܡ����|�M���hj	S��SRJ���zGV̦�v$�M^i��%~S��n]wx�h[��v�Qd�-�+�`��Y1Z
ZT)q<����<[Qw�n��9ZN�����¯��mFz
g�CjV�I�Hw֑���s[oA���uJ���L�<�%���[��7}�;�Y+���^�6"d�����mr��Ց��I
���Ǹ��7�J.�!j.�3FƆIc!�m :���?	whv^�y�y\gW����ʣm���Z��r|r�����ZhT��Q�]c�	EQ0��P��A�����60Bh��F�9�L���
�z�آT� c�;_�c��
]5Mh7R`:Q#E_Y+�ý� r��/9�sܡ|R���?�I �Z�%�<s�S�h�vdbR5w���gzJ�w��k��ۅ��E�����m2�B��ci �f��������mV2��:�k�ǭw�I����X˩�~��ƶ�p	���H��+��Р]:��E�rK�.�������,�e�U�$NXl`@��FE���#u&&��7y"FЯxN�Y�}ݼ\�����s,qyAAl���sϠ�dĥԻF�*+��4�T����.����$��T�����E�҅'��dˆ��NJ*�5�p�#�L&�'��M��;z]���)�t����Ɔ$�O6��3^<U���ze^r*� ��l�Z��fw��DwɊXQ�^O�5��Kc�%������������mAvೄ�"b��E��V�M�O��d����ǜ%�竎���J�Z\��s�O�?��k�0��_���o7
I9��&��ыw�7ݻb��e��� ���� �w�O�j�j�j"!|a�"�����~��F*��k��7��ex�,�1M~����IA�dq_�l���b��6�9��3�����E'mEq5@v�UOV����h0�)���a5㨽aw
-�C���S����n]�>X�M�b���l�N�
�Z��Om��B����\e ~tN'�ϱ�'o~y/�|P6�2�ھE,5����P>sE	����T7�-��i a`�m3Y:.�`���4r��L{��G���*qO"��K�K�Q�i�{����<9
�j:&�� a>%���]�Z�k����z[����$_����N� �� ��8l�S,����oA����ӻ�iͅ&�ɷ�H��$ב��O�g��n2����E�&�T�j4�X^[ݕ�YHgp����|�aL��"�D��:�F��6�R���,�â��Kܢ��HQ�z���#$��h���z	V_ݒ~�����]�H헚	�)�?~�{�O��||I�4Y:Q�1�5Z=�+�\�˳��H�ϝ�d����4Ƅ�]�Y�F�'~��'|`Q�_+S׌���֓��rf�ꬅ��-7�va7�}�{#FK��x�#��̇��D5t��D2�v�u����5���U��{���bA���m���}Djِ�=K�~�0�b�ڛa�	��\L��_Lc��moPX'���e�f?=LC�,���"L��+���D�n��@GgK}�C�0�����+�ؑ��Ct��d�*����}_�L��ػd3��W���F������r���t�]�������1���x͐ɍUj�+��K�n�������?��H�r\p5gŏ=�����-q'����Ė�{v�v���
�������E'~�<<�pɪ������`'�5ư���@�Ǥn��a��X�Vt!4A蚝��+��N4���Ө���8�%Du�I��ɋ;$��T�!)�D��w�U(@]Ǳ������.�ŗH��Ӡ&���2D�=J�7_�9 �VE����#�@��������IJ#�dz�@xfɸ����.]��I�0��萝Ե��&��ᓏM�{��uV^A��Ir��f�GJ�BCe��m	��m�����Zzް;�s��/[���7X� N�G�ƞ%S�=��N�Is4��I�*�9���#�CD�'���w�3�j�8�Wi�!+V�k�HM��ͭ`��^�i���@�g�]������n�D�W�ESdV���἗��J(/hmp��{{:F��w��`����G��\`���Y��C��k��]�.օ�c�y߯d�D�&���A�E��=�T�o7p�8�۬��.Rz�����y��*�s�#*���ˢ酿11ê�Aw
f<�c./�5v&��|W?�$��點gN�s�����Y��B����u��<�NZb��8v��Q���n9�񘋲�F����S�,+ҵ�a�K��;������]�*'y K�^`�&��G�s�n���Z9��h:x����bq��R�_l�|1��^�(�:�D� 2�u?�GX�݋1���^��D�X��,���Ĩ5���5r�r��pO ����������[+��Iy�C|����[r�E�s+�@���M����L��I�Z��x.�s(��@���\5a
���&�+}}|&a�%�.�e�@�o�� �<�	w9R���ɴ��Ea���<��lsv|������]/H�t���)�,�ep�m���F�z��3϶��ŉ3~C��	fj��<wk�S�p��O{���c{�����	�(\zf��c�Wk���U��
T���R��PWP��4r�hi6���%:���2�9��G:h�݂��y@.��T���~[��@Cq&UN� �`2ܝ�$ٽe�~ʂ5�~��FwJ�C(t��>����U4�����L凜N�4��X�үO�X��Bw`�Q�E#��Fmp�H���&�w�"�7h��o^��gidU��x��rF��#I�fu��2�{��IT�,j�ݣX\t$C����'A�7���^d_r�{Bױ|�:�`#���}�60�P�$'�&)�!���o��=b����=�-N���^��_MYz����V=�M5���@�d�̈�c��F@K��i��#p=�|&B�kF�#k��rr=�+#OJ��z����,}S�8��1��J����0�R�~�67@s� B�Q�6�VU�"z���f��`d጑n/4@�V���JM�u�$�����$��Ԭq6�z�m��_�YJ.oF�������T�.A�v��R�3y#�g��{��I�"�&[2� `��-$ݣ�pYv��"�j'>��GV[{3-�k7��#ZY��QU���~^���U|�D����8g���ߌw�����ҎC��Ō���L�^S�	��`���֦�8�;�0�����H%\��ga?�)�짙��,$S\��I��o�02ʭ��g�f˄�Z!Z��u%�W����^"'	[fuoj�NT�[��ڕ�P]���"��Eж�|�<?ݝu��d�K
�8m���]���^T�FG˂���;�D�����x;��A�ـKrH�O�&R�E�7���q�����|։���h���'y����-��Z4�v-=�Z�̓���*�=��H����&��	�W���9��׌�A}�}	�c̻�9X8 �/��V��"֝����۾ˈ΍�M���r�!G�^O��"Mt#�"��W7�n)�����]d`8�^��S���d�q����N�q4q0�W��lBS��0�B�Y@���5}�ڭY1�H�U�*i�萬��6D"��}�W_��m���w�F���@��p~lD~�FfI����S1�49�G�I���E=������� �shJ_�(�