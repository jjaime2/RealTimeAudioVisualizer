��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E�ﻏ��Aގ�~ބq\�l�1�4QQB��t�
�_�㬃1Iw�$�=�\�:�}Օqգ�$�ZB�h��NS%`2#r�e��c��B��FJ�CH"!��G�D�}��za�����<vri���Q-	�d�!�s��'�*�bOL qls	��{UŚ<R1l̬9��)��P)ۇR�	��� ���n�5p;D"���mZI�6gT��z�6�WLg45��sͼ׬��*�u���S�!kj/��v�!h̓v�ӣ���?W2w�1��i��B�ћ�����fñ�uCnԯ��&�z���)�?p�e�9F�����x���K�>����g��?�L����&�"���z]�%�;�9w�;\��|.E���z;�E���!;���+���i,������է�H"G����R#~+7E&���,HɄp��w�-5Cy�C�ħ�f��\lR� �pt��]HdxM�{g�Wg�2 ��Y\�(���ȡ�*.��oٝ�L���b0�e��)`��T!Ar.��y�7�P｡�g=��8	�����x۳�������Rrn��.%�kdy�9�/4�٣�Z��|�D���Dr�o���=��"��r���h�( ����<�n��]��%mH4,�}�R��!=�{Ƌ"aJ / �0��<1��:�K�:�^E�BpA�Х�>�C�;��ء�b�ݐ�-y3v�x�"�����d�<�>�9���1M{��r�?B-���V1%`%�TW5AcEu����G܂I#z�^1�7l����eٻ�GC$P���������*��_{�\^�j��+A\����c$yv55.qc��{_$������ON~��"F9��9����\�Ƅ4�k�5��~sC��W�>��l*v?�ڨ
��5J� n-�H���J)'*ј��6�q�]V��P��2B]!���^nϲb������UZ�p,3�����r��Hxx�u�R�pm��x�����Y�}���n?;
ڬ�����#Z0��t�{r�/_���E0��Eml�@Ey���8���otx�2���(>o~;�j�j�@�2��d��D��g�����e^"��ȳ9��Ό�b���@Vq!	����LR��m�8��I�O��V!�꽾BO@��4�X�?�����ę$ε�OO���E��R�������Q���|і0/��㓨�D������� �X�	�ĵ��2 @���w�q'��S^����(��L�����ED/��ј��`��"� �X��ʑZ�>���cT �Sנ���i!��� ����V��� e��.L�w��U}�W�!��T�F/_:��R:�@�]$�. ���H��	S�.1����,���������I��L����Zb~�guR0�e6)ȽioAfKV�rrL�qB�8lg�{�	��������'U�O���AW�U�)Ɔ�vr`}W�b�-I����I��<�X��r��sE�#���c�r����O��܍VӯI3���m��C!�PE�������B���-�o�:A�\r7�΀�qַ�G���._jj5؊�Z���G�ឡh���B^P^�j�L<D1K�߂Jz�0%W��aw�n�y��4_���a	[;u��L��)9�wY��g(��D��3�Wn֗��q��H;�6i�-a��#�U;$i �7rZ�AI]J�� z�͕>\&�|N�@D�|���	釆�D	Kc̒�u�'����X�yN�N��T����� :Á]��ҵ"���mQ#~6���8��E��7����ހ	^-�B�'�\Ԇ��Q�(�f�-6@�F�k]�5����l�λ��O؞q晅����2o��dQ$����he�cݿ�/�Y�Ǚ�K�F�dA�0��o0�7��&�������&���MIũp[Ё�(���������3�$/�S��W�r�zBJbD��_%��1��1(3Q�?ꁊW��cA��T+떄��$)��ϷD��M�����+�"�K���׏�r�"��84aӟFJ)$��j���Z�k�<Sm$�O09/��)�5��Y�t� ��'A3e���_֟�C�5u�L��N�uY�FQج�ʜcH�.S�X���P��c��A��
�Q��R�sd�l�.`���}�*E��&W'�Γ�xf�e���Bu�#q��g���Tg�`P�cv(1���P6r�q��i�;ؓ�?�cd���z�(�|��g�X�p_�Q2{0j�WHG�_o���s�5:���c�@
�c�D�Mh��9h�F�Cr{���ԗ��Jҹ$�0��\u�F�� �rm֦�o]���䋵���	�jD�ev��ڨ���S���М�N�2l�����@:��J�#�k:��⺸��Gl��<�]�I5U��VI��MC�%�z��.�K��
���-i��$���(���H�N�I��M����b�zy�!뗳�ZO�.h�5X~s#���Zj�Ҽ�(��D�r`{ð���KHV�m������$���=���Dv�њ/�cCF����c�?�F��(7��
�P�tA��B��r�QB$\�LX,�,c��t�Ǟ�3�{�!]#k����'��[o	*�ɢJ���_�mȶ񛇰�(Xc�G
	&X�7|ɀˎ�٨��@(�t?z0k��=�?��L*R�4�۹�^;>o{�+��@��s��	%R�a���=R���P���2�[׾��"���/�cN�w��
T�(]�+ő�ڇO|��B�9��kB \�p�@$�.�{*�eSBk���Rv�~0��ɋӠ�o%s����������#I�:�a�[���{0���..��~�s��H�z� _(�?{���3�3^��p�����BF�?�%̒9�Hs�I���L�U��d�����h���&1b_�׉�*Qr����h�)�tz!y7<�]K���}�t�nḩL��ͅ�m���u�*�SL^̑�R��xJ`SS��G��c�J�p������%���2��Ers%u�Tʯ��V����XN%����h>�{	3���k���ۈ���c !B�.�B@�5�_sv�x�@�Ω'
���K�LJ<�����0�l���|p�\6��)��!B|�L�9aCP���_��Od��"V3%���88�ߋ�8MR%&;����V��@Xx��)W������0���o]>��c��8��i�6)_a�V��\�y�֣(;�c݀��Ŭ�¿�j<X��Z�������K�n�O�7�N���7M1���K�fU��+Z�0j��}Do`��-�N�^n�=��WK��u#쐗y��E��P��Q[&�Ɔ��TR�ĒivZk=��
���?�V��Oq%A��]������9Q�!eR�T��
6|���#��J9�D���O����W�D�d !	-�1����|�w�Eh5#>���s)H�q�H��.�z�G��~��S��f�vh8ă��a0���>���M������ټS��o�e8EȹAj�5��������f��,B5)0N-�i�雫E��"��CW檅��uQ�I��5 o����g �X��@�8��n�|R�A�6,-��X�Bf#�O�H�.C�_|I�!�)Q.z�.d�J�S������#F�r�
�x;[��=����y$��ga��~v1=�A�����O��7�dD;��+�#��;���+_�u_�3�:8+���v}�y�bc9�FQa��|�t��^l2jb*������Ez�I�&�"�k��
w�ؿ=Mwn&Szv�Iu4$_4��y&����7����P�CT�)��%�`�����3,�3p�F7��G�F�b3>��S��H�dܐ|_��~�|
�� _�^8�ܻɇ;�ޯ�J
�2�jZr��EA� ů��eŪ�b�:�|`4��ƈ�$1x�d`���>�夥[=�a�b/Ŭ���#�{9Dły0|Y����)-N�*(���~}Wu�4�k*n��U�*7w9&����N��Z��������pw1�E�pY�ｐs=����	�Ѥ���N>m7*+?�s���5��Zt���"�Ζ���Fj����T_04�:O����������������iÙ���N\��7 ��U������ު�c>�x���3=�:��?���!�N��O/���G�#p7�pd�a�N��X�=
���,8��ԃ�~@ʱ=�c����ar�N���h��8���l0ʓt�#�~�~Jf�X\�>!7�����i>��	D^��~d�]D� 6P�	��6�W��կ �(���?r
���E|���y�
4ѫ�����x�.e>m?�p����ն�v����9�(��[�KRtY&����U�����~qNb��o��$���#-�PH�(:�"2����3A�L��r�ne���]2�C���P�{�e��H ��+<7�	~�*��#9�<�Ӹ�3:�����J�*�7�X� l�{ �(��^�3�
�$�&lٖ1ÙĮ�]�TL�QV9��*#�|����5u�K
QxP��\d]�/�}��`r20Uܰa0�M�g]݅*6���G��`c�����Ι� I~�"&1�Ĵ��^o�\e��H��ںd4T�N�֠�R����<ƚ!F �ֻ�#���Cc519z��i����y���/��|����k�_V��t�?�!�i��0Nh�O��7��N`dͅk�in��IN��W���}J�κ[��	%���#���U�Cz?����-@�^b��l2��I���Ur��&]1��}C�W���Z�/�iC��2v�z��B��5�u�m�c/G��!���f}^��&���y~:A��U���r�7��?��a�CC�I��Ž[��>F�ܘ�r4O��+>J����]��_ᘐ0��^ۭwb��4���OrbX�M�_�Q����K��4Ӻ�XQ���F.dwf�gO���s]�� ���@y��(�crj�~���\X�X�I���1ˏ}� a5 �wjL~S[���M�����V\�o���;��X�Hz� 7v%��p>Y�e��8����F���pE�7\;�[3{\,�R��s	H�o�����A�<���+��B؅E�^3z�BHlM
���ӽ�%���W�P�ߒCXP�=×�T��Q�����h�(hs����t��}H!2��(�\������o�m��'�y����OA`a��6��&>��(�p2�+�d%�����M]nX�M��@�{xc��7���l�Pd#Vc�{��i0����uʵ�Fҭ���aߵO�kS�t-���I��J���U��ǩ���υZ�(";���I]Di��w���Ol���]>]�J�^��y= w�2�[�e���[����*7;�})J�:'�^䔩�X'�ܹ����P@�N�J��ٌ�����}�\����Z�ϝZ���c�ݴ��ڋ�����&�6�Ē���������JYw��Ra�l���2��[̰���ş_�eĀq�	���]��_���:�8���B.�?�l��ǃ7�2`���Wi2���}��yh�t��U��!ⲥ�Q��<Rs�H�~���#!��N��"�)�Xj�h�E�Ƕ�[��^��$	�_nZ�E:��J�i��{"��~�	�a/M�JZ[7�|ۇf�QdM"yP�y'~Q��a��a%Y�{KO	��Ɗ���`�t�CV��o�o�<�j���)�Ԑx	��~7K�����15`��U�x���c�zO˪?'����\&х0Xi�|J���JM�����kY8��Z� ivb�3�2<�Y��F*�
��zc����F+]-���M������v/t�g=a�:>�kH���4� l��?ώэ��a�Ƹg�.vޒ*�ς"�r[ 1K�0u����<��P���9�(5��7�ݛL��$�;?�{��qVұ�li��d��S�+��w�D�0�1[��۫�9��!7fc��˟��4
�v����1���SkO/��ёj������.~��zC_�K(_I�����*F��EC�f� ������ݠ&��M��o�p���/>�Q�8�8�y��Ew䌝���$�ϔ��]];Q.t����a�qΠX�La|�b��,��Y��;+����B����X��!���6�]r��t͇e�yZ�
�9C��g�X�['\�	׉oS���G[�D�u�`4�ͫwW�тY�=S�f���?J�M,��!cf�}����j)S�Ar�����堡�yo��C!����F� u;H�7Ȱ�qMi�d�VgR���+�o�D����Ta��{2LtN\���Մ4�Z��ؠ�!��"Ȁ,+㤒|ʊ�j/ǫx��*V�ߺ=L�&� ~�r��_4cd�����Y	sX'-�u[|7�&ّ
|���57{���f�o��t�� w�۔+N�Z-�[q�+w:�;;���-|��� ��d[k)�U���P�G�_��/��aU�9Z2��Q�|,��
���뫊��FL$G�����4�a �^�C����� �����p��W1}p$�@d���S^*�&J�F|�5�vޓ��L$�EַW�/z��(7e!�Ό�x�>�Өnw�h����e3L����2���F�8�g�c�+	�(������:�m8���lH9+M�s�H�'�?̼.Cg��ߌ��G���;��_y<�i�8�֐"��� �H,�r����m��,Na"���a�?Gg��vm	�*,
$�=����U�o��}:�B[H�Y���x�~�
~^o���)_���K�Г5+����������(]�W�ԕƹ��0q0�"�+م{����=T��o.'�z��F��vﰛ�s�3&�Z�]� m�i|�|�]G,��@����h�ŉ�M���VBu_k�,5!4��C�2��+�|��P7쮡�~G�ޟ���w����B�,��xf��C	��2����42J����o01v�s��&=+�()ɤW<$�A֘�2K�s�J'��'�����Ȇ�+�48B9�+�R��4���젻��Vפ9�duZW�?�Y.��B�xr�TD��vY�4��,�]A z���S>lT���5�X|`���}���`T�U�y��I��[��W�8��-B�	d�AR$����)K/F�O���p!s>��ZC��L
l����H�%�s�?�n4y���2� �=-^)o���g��c��]~Q��Z&�;�mR�x2쒟��	i�fM�wD�R���G�M����)!}��k�>I���k�6�AAPe���l�6�>sT����=Qx��Bc�����B��Xd�>:/�sn��&��(� �i�!�0���t�*�P��_@.��'lN���.� ���CCeX���r�����P�d ��VHX����;w��ً�5�;�y�s<��o�Ԡ�=S�#���<����,��;x�ܘ0Í���/�4�g�B���?�e%q��� �Щ�ڍ��涛�s
j~�SHK1�O����v������l�ЩFt�G�R���k���A!z�w�Ǝ����d�xP�q��Y���g^4�o��L���׈�6��
p��`��5�@9��c���|�ᙩRұ�o89�I!��ݓ�O��ػ��|��@ZƉ�u�99����&L:�pؑ鲜Z*qɎ}L�m�sR(�0/ՑHg�wA^��˨G���Z�,����r�(������/��#qv�v�Y���/m�J�:����[�{?��������RT���ⓡ`��^�в�Y�4.8R%t�H��8��EwZ�~0��Tx�s���Q���b@��IoN��^&�L`�j(��/%vy�^ǉ��s>��c̓�?m{yWU�;��/�?P���5k�⦱���	�Ԍ!��U��F�R�+��0���f~����#���}���"��ޞ!�$*{�