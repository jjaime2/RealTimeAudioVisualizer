��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊��5b��rt58f6���;m��#R��pIKU����A�b�@��N�6�ܲ����d����^O��	Rҕh�|�4�l�MG: �8����<�֯���~�mK[=�)��N�.�t��]oannƀ�!yhu����@s&�P?����!����Md�wo�}-es_vă1�h^�������|���I��hD�N��B^�@}ɪ��3竎�$�*ݦ���ucS��N��8|.0~��Dƍ�/�礘�FeM�3�UoUܓ�����?Q=�3�0�m��r��~	������9ևJ�̸ʛ�V�%��3�ɇ������
ꌮ�wq6F%Kr��l9mqf�2�&�W�[��[煀!;pm�ϙsϗґ�UpbJ���K�j_��}��ڎI��w����˞m�!׾��E(䨦p$�5-�i��\+a�&[�s��"}�A�5�Lcr��"0w�	���Û�����O���j�b[F�����J �X��ۂs5���U���<^�@�0���y��,�Hʵ��[0=�d�(�-#9'�&�������jYS����3�?4�p�K�|KHj\�;�S�Ȍ;=���xZ�Dt���4���Zp[ӆh*�������:��'�^��VK�T�K�@W����ODc��v�u��w%N��H4M~6R+�7�<�]�WCh�&��{�rVK(�f\g�:$�������3s,3�ge#��_�7��%���v��ԕrԯ��<��+ԸN�C�pp�=��lbE!$h�{�ͷt�>a�����F��;�H�U�%�|+���_�"�V��G�R

u�9�/O�k�&�%Y�@�.��rVFh���_��fy�d��*1,({�YL�2�x��诪��{w�{����m�����?!5z�UI���٢`x�<j1�}]sXye��ڜ�t��3��E ��tGϹ&�!-K��o���m������z~88c�z߉���oqn����zY�����;	Pi��G��KY9��c�1�p��I+�8F�|��*�z�]��!q�+�j0�f�/��+��`?���n̲W�H�AC�dZy!��Qu4�3v8DMb��꺨������9x.Q0����:���S�:r;}0���9^�y�J7#n�8����̯3T�Ĵ�)=c 0	.�g1Y�t?#�����]}�֤��#��#�#0�i<ޗ�4�1Q�1�M�g&g�
4�V?�K��X+kVw���!��`4Rx�y�֋&�U���������*w`n�Ol,RQ��)�[h���|4W} �"�B��V��+εE��jj�ge�Y�U�rD���1"P�F�Bn�ȀM��X�͎�� ��;�ʂL7�*���ϞC�K�x���|���-5 FA�0d9fe��ݨ�h�y��J�O� �.����2���nAG��ģ�<���� 8���yᕥ]e��`L]���:ףm@��{��������w#�G5���Pi�X��.&h���/����K���*yD+�hѴosK���~���M���#q4!�I��")�D�{�P���,u9��i:�C�]����A�2u��qO�O	�a2ͤ�pmKy�	zx[��AN��"ʟ�j��܄��t�ݓ|���h�	�[G�o�4�ȁ;���$��;�i��ǒ,ĸD� X\$����N�r��3;�sL o�ll��(�Q�%){�@Mxɡ)m`TU�=���U}����o�  g��I�Y���$P-kIܙ�a���hUZ��͆m˒����JG�����xGf��LxF5>-M��
^�D��=z��я�C>�� �� %�; i��#�P鬄��1�3�YF�3|	G��B(�����_i�Ջ,&n����N��צ"q���3_�S��TNTW��߳~�@�!�꧷^��"���yk$��5��Et���+; ,����nQ�)�Xȶ�Y8u9��U��7�0E�V�TJB[�2�Y*�#2�$��x�"��"���������E6�sM��X)�/�~�\���B,3���{,�8@��	���w�_⃲�g��*����:�F�Pr
�І%)�K��*�siJ�zJ� O�n��R?SxR�z��\���@�YN
��8�r{��,j+�Z�j�O��ݕ��ͭ�~���a�#��櫉
���G�Xq�G�=A(�笝r��t�nE�؞
�?|!�'rr��i���{��݁q�����|���^�����T��o�e���Ҽy��R���o�p�,�F�tėemI=k�,�ZHyR�D9u�#��q�P�6� w�ow��ۥ�M'q댣=�G�����Hoa@��l��XbJ&�M`��΁��OMw e�����(^�-�Ł�C͖� �"�M��7�D�k���KJH]�V����DS?2^iP�)�׳Ƃ�1E��`�h��x������k�����\�5.�s����� -������\�3�����h"`�~�|�䟘��d�O�T�bǟ���V[aS��3��� }���~��+w)Շ���n�F	��l�P���=�S4��cۅH�|�H�E�����?�d�+�ZL��*n�f�87����p-J���dT<����b|{�:�/*K��gȊ@(a�$g�&��KT�d����=�֧�ª�B��!t�\��a;������lUeU��D`�{α\颫�ܟ�!����r��i�����\�k:�j����n�t��Y���x�)'���\w�]ر��*iν�{]�����	��#�aS�����דX9��V� �My��m?�T�E oG0�-�9����U� FcY_�|9Ҁ������-�ɂǁR��+����Z_&�|?���������v�8�@�
\N��G�;Y���E���GY[B�PW�[��7�����&��`�;�*3Y��B��w�Ȫ�q�o���jP6��E�O|b͗@���V�}x�%7n��"&2�f W�Q��*J:�G�O.�C�%��aY��Z�D�Lr,���zUǠJ._�KmZ�����T�x衫w�T1���By'y{{5X'�2��hc�cyG]�_�,<p��:��e�g��z���]�c�%%>S�����L�c��a�f2'g �D]�̈́cD(�⼕�qw�f������a�����H�k��s-�4�+��g
��=ԗ��蟘��V���E8���N��//���rq?�����C�e�(;$o�+�c(3}P���s����ECP�~	﹵�z��[vQ#;��pvr=�cMU�7�Qf��Cd�D���h��a��e��t��L�dy����r�dm^����<�DRs���$Ο�v}��f����_53?#[��@�tRDs��m�FCb~��9#�<�pW8����`~>�n�+���u>
rj4�Ii}��Z&֛q��5�`y8G��q�z�OG������^�쬭�xմ�ڹ,_�0�巌)��y�m'\Hn"eһ�[�:I��IK��0'����
 q�^Z?��5;H�D4�;^2�����
=O���ekJ�e�|!j<t �hWP�ѡ��1xKx�IaY�J�:�ma���:�������tܼ�^)�7'�S�[��FT��>JK���J�^[���N�	b:sZ�"� `cu�$��-��2�S�u<�^�S�txʌ��<X��J5{R��BX���pK���/w�A0Y7�����Y4t������3��O�Q��/��.N�_2���.qO��C���<�K[n2��&M���`�*�~�H(j|
˙fp�ˑb+��E�rO_\@���c�"
|��d���Q��2	�Ood���d9������7΋�h���_��]�����C1X ��BZ�mda����b|�"v���dS�%Kҥ8�������'��%7#�e�t�j��Af����f<&۶@9�bRj�z�� �ٝ��
/�������RÊ�6���}��:qR; ��gKB�o�.�@H��!�_�O'�c�#̬��!�8����Ԍ^�ʐ㫰e�(��-�����։�i�}(za���W-�X���Зў�����aK֐ݚ''�^/��* ����� �?�+c�cpH�u�|z���m"�W-0Z�~��_L�%MBK?������B�4'��4*��qϟ@��Rg����^������׫|q#�ҩL\�m������wt���l����x&B�GAU%AUc�)��GGp�K�*�_��%{ۛ�X�=S��Ѹ�tT�K֎km< ��P���۾�ݳL�l-�uQ���#���eO��/�h�S�cC�_"�.{D���T�K�j؛�s�;ꟙ3���˒�@Z^��xʰy��<��g:o��{��� 8[a��l��!z2�9����Q�6��ݕ���J���S�н�9^d�np�#�$WL�S����H�Ec&�-�*B	^&B�O+����n��>ܶ=����u%��h���$w�URo�\��N�VX��l����ػ�'c~i�ܛ%�����~��f
�ӂ�,�n"�
���2Rf��;7#!��Kj-2����C�����U�m�R���r�fq�ĚzfX�)Nv��k�6:��P�ʩ�l��:Y9<����Km'W*��l ��ܽA���# ��˲�u��	��ʠ��3t2+{ۛ���,A�A4���y�)�n����(b��\Hlp9����~�_�ht�2O߮ݬ�T��Eգ�cˮ��B	��։��,U��]�)��S	B��`����X�Hõ��6������~쁕>�,��5S��.,P�h�����"Ӛ\}v#*���/�8���b����a7��+xw\$,��f�f鄮�uQ�p�G�.�RUJ�h�N��75��<ƻҜ����y���d�0�K���^��/17z���Ĭ�?�);�q_����v�N�uU�b:�|��h����^�۠����}頽O��r������E�����5]���֝;���@3�������<���3Ū|�Qj�-���Fƫ��)���0:�G[S?�'�.Z�Gr�~���G|���~,?QfƩ���Y�S���N�X,G��^��+�躹���<_�!	~�M|r�+��ù��xVU15H�Қ�^b���ԯMD�n�	�.�ٺBOvh��m����"�B,�8�ş��D}�$r�;
��A��φ;jej5;���E����=��O���C�'W�YzL�cR[ΩEyF`TJ�Ǡ�WA�J�sf?��j���}l�g4L�O!99�5\��˞�e/a����y9RW�U�^�K�<)w�NL��s�
NP�}�Т�*�Q|�Uo���O4�"ʤ��Q�)X��o��ݎ�m���\#IYPY�(�T�������$��!4<������'WpS
�>��ǅ�T+�T	�I�Z�N�+"�:��^R�C�x5�|�[���}�RG��_C��Ǟ�y]qXט�8(n!��'�s<U	Nh�H4�&�k�����
�"������cԀ�VJ/@~���\ҍ�P��+f����)�?&Ht"c2j��;��17uw���`ֱ��\z�Z��j�à[��i�ȴ��\�t�S�䎹����d���
���q���m_^���F6���@ƨ�+���R:*�<Y�NkbGi��K��H���syќ�I�Q�*`W�Z���9R��VC��^�ɓH�q��DX���/ 	ZvDr�j�õ7���퀚ٶic|k��p,���j�{�g�,�m|���]�m�ǌ�QB�R��4�JBa4%�s,��}���s]�n���I�=�l�h��v�Oe'��e*��%��QW��W��`�q{/%"��	V��`�q��NH�Y�ŔzS�q����e�T��zy�Y;�?�cw��0�b$���ڀ�T�l�Dl4^
9bH}�P@��8�z
%�^��&�"�4G�C�W��!Aetd����%˸.�7��[M'�EɍX��U� �(��R��JVj�������,L���E�fzn.ڰ�v��$.sa�/D���E�-ɛ~YV���̞�?	��HR}���Y���^ƛA03��� �ې`!G��}m���@��&�v�bAO�J�f�,��V�K�5�[a�g7g�e����@�Q��	j��m�଺4ўp���j���O�F��g���,\SB�ys9�Ҋ��Z�&׬�Ve
V����_ ����ä��i�:W���c�ܧ楍�m"&�CJ��c�m>ɟ�&�������y�����ǥ���Hz1�b �������Hy��R�F��Y�>�Hn8	�*¥�xw�f��7}/A�����WX��8�m<��:,�ρ$f��
s:��=����/�}K/G�:ŉ�0
]z�d�1��nII�Z-u�Pwf���)��k����p���Nl똜��q�8�n�>��J��S���Nx~)[E�;ZH�3Q&�$1�w�0C`"�D�<u�``rjP:�B�p�8�=��,���?|!����k�����{��Tcá�,D�W��u�a0�-��*a�E'!��ETS	Q^>��](�!j��Z���5HL�,��ْa���5��\D���v���)�pI��A�Y�ؿ�E�;6��W�z
2;Y'���ǿ:�r6�j�<C�惏��Ź� �=8n!I�M	]��#��%�̆�����5��t�T�ҹ�Ҳ�<��̤�rO�8Z�w􎽲�j ���Ì(��v����g`X1�w�)��ƀO���=P�=��]��� y)���G��e���J�y��si;{WV�Q)����P�rJܨ>�J�C:���:@�A]���'�p)) `��A����s5�j�����q�Īj
�F�T"���x�XT��*���t�8����_t�X(2}�(WL'���,!,n�k�b���G�e69�{"�_a��]��YTu�_��b�E�غb�?l�L0�+(���h���g��U���j�"�g^������L��W�
S��Y�b�˕�ǝu���X���sc�X���7;���h���e|6��R@5-�R���8�[��`,9��\��p_����]������w&������H���*@RR�n�3�����xx҆'�������H5iQ��B��Ϥ��r�iصf�r�E��
sjf�ދ�B��̺��֖�!���
�(�0i����+�OG�����\'W�6�gVs���,�����Q���c��[�� K<��E�P�^Dܽ����n(���0��g^h�8;��$�:(3���s:v�9dhJ��u����3� ,q��2J�%�ȍ��>��,t�:^��R���1��BM����˫}���b6�g�B@L�@>��������8�p��1����lN��������tV�"��pԔ��Ǣ�P�4�a�R}a|����|9s[gY���_q�<s��_��m!Q*��3���Y�8��"0+�}����H�ج��<*>��r�X���{!i�.%��P=L.�A4�t���q�������"ޖ���y�􁰄���������������sS���� Oām����Y��ue�Hvu�J�u �ӹT��JBG[��0_]����ѝ�Ae]b�w�]y2�Q�T�^_��tXy��i� ��l;E#|a�5M�-F9�qU���x��p{�ߨů�gNp��fJg�P���_�o��OL��lluR�,#�F�N�|u���>1�L�8��)��ֆ�5��CI���"�����k����\��&�ـQATzrޔ�g bH0���|�&_�i�{!�1�"~"�y4>�d0��S�Y�섈���&T�BV=���B@�QN��e?w�Bd�j���G��&0��� �f��N*��x�Z��� ���`pm�칁C��@�!/_�����s7�|��5���`��	����v��ԑiQ�V`�
 j�ef
�nG����)�Ǹ��a7Z�m��^��:�qfS�Zo��ʺh1�'�%)��B���N¶��F�<o�s�$�i��O�é��r����28&�^Ek��f^���nH�g��rQ�yϕ�Փ��jE!��D<؞D
5�&-.�M�o��c*����el��m!��.�l�@���0*[��A������z0� q�c=3��+�?&j�����S�8:&χ�j�g��okť� �W����W����:��
b�I����uN��)ryr�.,�Mrk��=���MEY�L�\\Q��nA�x�;��۱@.મ-@4M{��ږlo��ı���Rm�
e��W��@�KK������'�Y�1%�A�%�$��94.�@�W3�4�n����?�L�3�_]I��'�_���%�'*�4WuKS㒇�ϔ>�;�\S��y�~�l�@6M��P{�N�H�G*�iUeвi�!6|������@�*�"ش�G����V@؜&7�%Dx�0��ۆ-��"��(@N`�a8唗��ʌ�f$��I!�2��/nf��[k��P�T�#pY/or(Ο����z
X@��J4��,e�Uc�Ws"z���n���L�e��� �o1���l��/�� ?�d���E�RG�wF!��m������"&��#Ӆ�	Nq$�H��j��g�K�e����X9b��hcG�a\|P�+����/����l�=S���ݎ�}�m�>d�k[J�,',,�uf�j���3~}"����y�6:�ʦ#2t�>YQp�D��f7�;��?��'	L� ��V]q��)��G�'AD�ۣ�!!���uI��4rI��`i�؍*b8�$Lh/��|\(�+8��l��2�77Q�F�*0��
�'���^�k�jD2��W6�"�ɽ/{�p�]hr�`x����Ҙ�`K�NI���Nݺ[���V'�:�H�I�	�5,eվ��Ͼ�'`f/[M�k�������OYe�:�K�l���;[w�UFn���aE�A���8��-�w;�%VS�����#�w����(�~:h�X?oPǻ�������v��cRa b��K�cgiSS)#��R ���5���E�V�b��a �3��z�KЬ���w�%� 4��H���i��Q�ڿ/z����)7|?�-�eL�i������w�j���r�v+-h�=���yԛ6WI�#�^ ��Z��⪹��L�Ӥ^���,^�BX_�騸�yK�;��9����j���9��t@�C�����"�V�L��J�Z�ߵ��e�Te��͌v��y�nX�����<$���h�/��2�o��.7�� ��C�&�;-6_�m�c����q��q�L}s~>}Ln���Hw���ɀ*v$O	'En�1G�����
 ��&��
�x	C~�L!���f{�r+y�*���y���L��%���M87%�18���}���9��OWwmF�(A4�	���5�*�Eu ��kK:�[���V��/[�SѨpm���{ƹ����E� ��x4賦-�;Ǯ�
[t�"
F���ND��Y�-B,��p>5(��Dm�x�������n�`���{�ʷ2O:t����<��n��w��h#�HR�������Ȭ��)u,�ـsF	[���.$��o�h�L���:1���y�c�Pc�C]�I^�RC�#5���E��H'�/`������-�����>7>ŽQ�%���YC9ӧ�N�ͻ۝�7��P�a2��6m���KR� ��K:�G���b��<�O�k��z�.�O�._��kiI'3:������Q\���=F�i����әl"W�	�Ѻ�X���,�ky�t#)�P)`f��������r+d�y���??����PH�s] 	�.W�! ߞ�Sv��+��1��n�B���&�����IS�V�݇���"�(���3��e��m�'yO�<B1*�[�UWЗ�j�X"^?���M���h3N�ގn������1J�ݐiyB�a�'��/�0��7�Cm4Ak5�����.��)ƶ��$��[XV�8�6OV/w�vߚ*Hyz��D���O��W�ЎԿ�����-�Lv������[���`-�
&�c|n�~���H��(�׹J�M�ޞ�P����...a�k-F�uFOB�)��@i��(��h]N�����q_ �/Ht�����@U�Y%�z+�p������m����:d0Ax�/��`T�ֽ1"qNng	�:�	(Ƿ�ԅ���|��)��`l5�d&L��q(�����{��N��ڦ�Eh��.�"��������,�c��	��~\k�%� �>