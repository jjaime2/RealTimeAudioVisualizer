-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LDnmy9pMFgCN8nnz9jjd0tUsv0CJcZqXdr9LI4/Kd9eZmF0eStsJp2JMHY6VhxdN2WQB7d2h14hf
9dHoKlfmqHZtxGmss58jDTWEzPKxzhqjFQP4Cs4sKsTnBgBBX+0KNaHyRn3NBgZcCMIHa1O6Ete0
8OEltzAFNRioyDsgnODWpcK0mwl6vCJ8GPUoOG2dDY6qdRkk8+BRPFlgcLdHEbrpljrv95ywxPOn
miwR7VpU7rGTz+ggrIjk1UrB+4Y0R95utcbIM68vLfvAHHzUpPxKUuvgAlNVrMoAUV4FgIMZ9h36
N3mM+7eR2QIN6xqV84gVL12UkQqrD8rBXEl+ow==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 22000)
`protect data_block
DXh7z6VzZqsJYjtpPl/g/iyHi56tSe8xss3JYh1Mv1vSqq0lXekLL8TW5fMeglznCjdmiNjAJYki
UzCLIgWjweNJE62FJAcvL5QRdeaHqwCm4NYzAryRzXPHiSXPAgQqE0W1KZ/WhaGaF1QoqN1zNwSt
RNmMmk1uaRvvN8rM+v5FqvUiZj8nhIzAMGfL7LAZTHP8kUpXMdSa2GTOoXD/Jmp9/U3T6YhGf5Mh
LdcoMQt7HQYYBdK/blfndJqQD7a+sf/MWMDwVqSGsrD1cqlPiTQVnmgY0R1hRHRo8VFlBWm1yEVH
rKByRo2WsNzj0bzI8RCHFc3gDynsirLq8gXI1WOunG+FFuBmM2SeLN8Pb9LUxwJtTL6Yr9qlp5bM
hIraJgejJa2NBArKjoJ7wQd3agEeR8ICTcybhhIIcxzcerGaV48YHGPhuo12knwr3SkguQKoOjzy
OkxQMmGJ4VQeT+c1cYoNrtTm5uRJfxlN1J/yMEMzIhBWQPYRIqjqzf/A2JoW/vyWp2Ld6fAl01tv
pj7BaZqB1bcbJ/K514GTWjPvlNcH2DWmGDqhADiz2NAhK+Ox6pf++nLhpU5uhVdxlZXiPYKeS7Yh
j+Ha3VLT0RKXW9ZWQEKyOJ9LSshZgnFjP9i6QzgFVe9Z6khDCaI2R16OdIFKYnWVKEFKgIMx7rLc
2NEhKeGu4ZYM5uPL3xR+xtmg9Y678Ac0vA8f0dEQ8GBSFgokN4aiCjtXNKskBPZtnSvZPitotMrX
I3kSBggtH+e/tIpuPELS1OG+/uziaaB97pzhJqAlWEQ0rcI9n07/6bzDpNU7tqnz9pkLaRAGjRNP
kr4bL1HQ7g4cuug5glKQUE9Gvn/NoiW2NRAu8kmLfvGIHKyUOzK7rAYUMaWWxhaCeneec1qRxM09
rUY8upTBNUoQAloFf8pa8y1Imb4F2XcyPom6X8lL28DUQhKojqbuzsub+2D71ImWsc+oCPcjttmz
ClZBD89t5OhF8euAQmul9kbzEplCbrx1BluQsybasF3FSDTcFGEPtb2RhKaCm5jNAiu4MF5xEg+G
6qtifscN7YLo6QUT3nyV06lkp0avfCeA7QN85JgBc1mmocL//GICJtxbgeCwZAplL8MzCuJRrukJ
wLOtSAgzjSoW1VWhUM6Ilnahyo/55Yx5JvEh9xxTG6t0AsWnOnFF21WcaoCaxX2Yz1mcNTineMbN
KSOaqyFTXI+yNp/XKrToYk27lAayK6i7XSS3VxLhmAJwWnbIYMrrLwyA8CKpWGmNrLQ1yHjcJoYw
xybg2JuAqJyRabA5F0L7Pz4AsLDAPziq+w0JUbJaw/F2wVatLPLgEOJvtfnBLdwkWfQE3S1REX9W
w1tdvYdgMSjDsTn+ZHY6LyZL5G1TA8plcwVKo2Cu+SlyVz/7Z9rm8MR8PoTbs0dXlip27dNwQikB
L3uoQkO808Xuk+o2vRL9UCQqU6Pd2OuPJhgrkMw9oGuobGUniDOUML4D7zEATaMvuk/7L6EhxA5L
tr1uX7XH80aA1oxd1sWm6y7+32ZplbgGCYg/0r9hgtpNJZD1AEv5IF/HhoYt05gKWqkQme6m0ivc
DPZNdAY2VZ737OA4Zb6t8v3R/ag6CmwZRi/eAee7fKR3xVTMA9sVf6TrLhhFrTy1d38JfaeHiyV9
sTig1SjapEcnGQ7uCYR2WAewnb7ZzFPzlCuh51xAU81002j6l7a4aCsLJxlDIsj1pvbBD5cc3N3D
0t9Pb13IebtkM6a4OlzXKGJJ5NIJF75dJ5yBCDwayZpEFaydCNvJxUORTfz43rVQlwJ6+OEGiXBW
LbYl8n1/SGx9LYdn1LQSOLG7AIKbTzUN7d4K4puIx+Z2+KPhOv2AY+X2ADyxgo8JIlV6NY4Epc/K
iPvU9kUNqGFssOoQzsCtHcH7o33aDnkX9KoEo+cHmGFads6EOk5ID4T7RwhbGwbwtUADhRzZdWwR
ZGgIflrTp1uBusE+X/Zy7KyRYqjK05n3ZV3keQbi972V1qWZywgyFV7Ykc479Aet/sUZ/ZVm2sQa
YLWFCm+3eYKFwCXw6poK4lqQ/l4CGxXGkgq3PAyvn1YQmQASzoPMsS3ptwaZF2+sIYKCalsP5gDd
wnoo97fJb+SrDi4WeXB3OcgbEYpextesEFBZi9L95qUG6seDt9Udj5MsPm8WIDuXTDFdQXeXijZ/
5P9yOtrf4nHwJecnwk3P4YAZEhKoVXOH6EEOzWyNp/w9wMUJSPvIbmLCfAlPBqLAQe0uGiE9DkHL
6d2dh7a5NACttt72Wi7z4few4hbvis5Kni9pgLRj1LDrZSjBaCDGHkg1JE2uC1x1MPrj1oN3F147
BCVEQ7m9piYZjLekHHR0pC66I3W06AdRb69/WJroQ4/4NijqmoNWAcTQwPydbgZAWUKWxbHORPK0
wrLwZZvsT+1PYY08wn3VFaDr7SBHpZdtTYddoJHv6YFf4moW8OFRtlGfgyiJoQvP3L7RJI9Ti0cY
TsJBD0UvYxl6UGfsTCFnz+g6HYOeQPTE1kwrvYheGHlo/DfWcklRbJUGQSLlQtw3HGWMJeTckCuB
5/fk68ohzSZAOkfy8Mn9fmvrZR+8u0BeHXSbZuT7FG5/OLsVX56fHWL7h1Rsh2JTk0JXTfvbd/YP
gSzQ1F5HpIgEbOnGRbra1Q5lG9MO+8eb/4XoZDNp9g60/F+jJgnHSPDQtNXUPESmVMDUPi7Hg5P7
r0tCtqPvZbtLPICcF5nUpVMBs3TnXR+jvWNdiI/eEyWPt2zHBFRA0ZSzsDKJCZy/32jWn3WLyUG0
Gr2ZH2muDKEM0S2qXzIQUAhcwnJwpI2hxoqmS5GfP6JAnzCd1OZTklYruQXaZo85wO+YSJNFblF8
a/bpieiHwC2/qZpWhB9VVRQb4hHWat0g7QUTUnl/J0oTIgBIXJpd01fsph8Ldd9zhjEmI1ixEGvG
xCy16gca8kuFYYZAsWmfx/0kSS+DfEZ4/7FVgjwSdwMHljkIs32QhCWv2/RRvSqgwbe2qp7xZfEF
nMBDF3HOfA66zk+06PbcIpB1QfcuAetfYIDMeo53spWkfnS76x5z6VMqkZgNqyMCZQCj/B9FyS8N
pTdWTA4DI43t+rbKimBrnFt/mLn9BzxsTc5527c00mor1e7gFZ7F4Wd0WuDSiMjVO+A5oXmYZTBm
rwoaIGzTAN779Uqa7q/EBxyxLnOrhAAbx9LrxnQSVohMWIIZV2jS1SrOA0ymQCxLtZdPPBApqGO0
8gnppdwi3dtcHWAfwGhXYaPiw1KBxatn3xRUumJiBrrKyhi9yyeFpytsziAUVQ5Su+/bqDSSyk0E
V2r9CUFMSvsOh3ISB+QXouYlQwtc1nh15Y1eQEEQBcNyxdQj8OurKNbCrRGH468/BFfRXshmtaA6
zWiLbTijIgmYK9Fae+SrEVI4jvP9Ej36HgBNVSCsQDQvQ9FYCOt+jFsM6xKXznfEFqsqNJqif5Pe
ri59K5KV+ic7D4aYra1cw+JuzL2E5f47r0fHiGNL0XqDtspOEkF8RF33rcfhHXC9ZbdH8aSUtd7K
t4r2lIxNeeNhheAFzhKuF8ivMJbsauq+2/0EVEfwV/Mycxwa0l7KKgzDKE8SwUb/DCF78bzU1Ydq
w1s5i8FfBgcePTL2KTt3hOyMgg4VBOX23wOVcj7qaA83RJ48n7FZUs7sUb+CA7tXm0YKvUtACgkI
BHlYU1HOVLiPhew7X8Q4Rm2eyL0meCe3Y4w9VR0JYVVg5l0heC6SoXmnCZfnXWGZac5QE5DZnTYa
Dj1gkP8ZCpfMXZDSg4iZiS0nZWuewjxbW61wWeDCKKJYY5wXZqWlwkmbMDhgof5ojnQhwrqQiEha
6gxSvdfp9rXhfyuH6TRFYVPh/0yrATjB5HclU3nnXoVevkGKMnw1CbGZVi/+ImPvo0sUDtX5ACGh
g1v/n7VAL3M5NYN9GOCScIoQpCFy65Ki51VS7TASStM+Aj4RRP+Aq9bGw16yKzu3K4xVcJBf5yf3
H9bMl+/qInf+QdEwcGmOIPFfbeTKhgSRcgFjVg8/o2WUG8jWVBUWU06kGxElnVuqQ5gjP1UWM2ew
e8AQHpA4Am4uDeP5IbPlIRgx5jiMHaEase93dX0ltCPwi1bFIapS/W5uL2kdB0CVOLgZtq5l+684
zxsBAsa6ra5Bez3KRZ/cGEi0IZEYDoFU4nvNy9u1ZhGSJwNQmFqt0CUPbh7vPcaxmfHho1oI8v2e
uxN0SEEYrBGiBCtAm2P0XuqKk4u4b0k0NVSvEfBPOfXYD8rmnlu3LbqkhrVWB2kmccuXA3iTF4bG
8jYY0vWqjTwctSouVoFGy/dj144Wa8sHYSnAB98AA9MYmoeBBeUtdfmxJuObWtFKtPP9AC1GZqCn
z1DkbKhvUAkLKWOkvWJVpVilhXx4iglMDIzz/PT8dwejukfTgBy4wuGXqg3VZqFdmNgVMBeR1ke0
mYnoZCwjma95do3AhQOsRzYYv9G1kWKtWIFR095vFPvMouZV0kTnHtmEEW0vzxbEmvEt+47abmFX
MFEF3t2xIXnlNC6ova9JfhSVvQHKiSpjZyQQlvxhL6eHOjsKBcf1ne2ntE/ZFGsRgKCAhYpNqGe0
S/wi39SN8iDxNDsoopyMw6A4jCYURlYKPeiY0Q2JFE4vxLuH5EKc1IYg2D4Q28d57TXD/ag4WcUk
KRa6d2Fd0zJ+/Ok0WThgLt7bZUdJGLdrrn1kG6hr+UQH7OVTauUIsoNvsvsMbU+l7ZV8BmHdPYA4
bX7nmVTHZ5jdVnsS3Qv2Nuxn+eBLjs125pmP/3hCnvYgELjtnYxwgryi83gJwxLnn74/gkPtxlPk
h5rmgYGSVHB/sZ1FHidtBErfY+XQcE/cDOzzGf4SIccI7a52Ys3ZSI4dRKM+kPyHJ+h11Do/lwdT
wDNbjMfQRnMU2nIFJRO0UuvnWSIfNy1XQWsY/nOt/exxBxRKhRPYeUHwELwEnY6RMl1zQZKg57gP
w7E5NsQF6abQpEkELWHZQtDHBIrUeAWk39qi0GGUe3D7U2Q0r7MXkt1+jNegUQjxvNYnaemxluZe
ZUihTRLMkHx8bNSCZkcBpWp7VbCrUWn2lTidjHzSY2cDKS/V+GR7xv/SVsJxPlM4Lj8lu+eNeMOI
MQPKIvwA+yyNYysnt6Ps4f7T0pRJOgLpyDnwE4D6Gt650TCqgWX6r2sRXOWRU4YbphvEG0YKrZiC
BqlNOz/WXGfvN+gBVvIPjd6g7Guq1JGGtuCup0pL9IfxlHXfGNQwH8MfndHDoxizDxIxAdKmumsX
TsVZbsdsnS6ZTd1bFVdhn5AIxM0/JkQa+x4t3oF2SOgvR4CQwAXayog2pIifEdSz0rgUrG+HOF8i
xGHWm38UblTL5osXVB/727Jmy8AzWvfm5UyDJ/y9VJ/whkOFyogN6GEs/Zn9BWeu7frcu0ASI305
pdH6AEu8S5td7WmjAWbBlioscVj4Gt+S2PZgNOC7xhL157QE7hREFdiJVbYbSTeNMXNnm+lJ0C4C
E+H38ykkdeVLfy5LDbb0P9ZkM0FB7zGYtZXSZRQZleVwy94uXSAqMpMmpmtl1q3mAfvxN7YtKFej
3i9Xa/qjV0Y6IQPhjpFj4DrC/5qW/WAvvY7eIZHWuN0YNA0HfcbGehguxKCO4Iv8Uw6xWGpI3hp7
bW2DK9p2p0o9ucjkWWYz3UzciwMU0KOD85kaWdNoyfdO61WWXvTCZ48Gt/K4ksWpb9n5oVZ7bJdN
nW1reqrfNeV7CHA2IxYJnurL82+6pAkCofNFmYWy7EmLJE0/lq3072yFjH1EGlO0txufRHgqdoll
31RQxk6nMbgai13Edo+YqpdcLbBMaOnshMLT32kNfSFh/SpjZG6eTeEGp+z3k/RESUHs3z6VoJYL
8Dh20W/ujEF+DYHPIeWGlVsZaBmNv29Ktkiz49X1PVLSaTkvffqGXwDS1G5BTWcfeR20dDEbeU0J
hiRcN3J4ru3LYhiGEZHGfB9vWt84CDmerPugLIDU+f+jIHd2qD3kwD5LxFUwviINCbnqdx8ELy0i
Sf7U9AGqMvYWVXiWqHV2Rq0NPIVneuVG4nEcj2d95oiO3tl6Aa0tnuK6V4HxTX2Nj3Q+NQ3mZ/pz
wF4FxDhrmFp6XeoHq7pOVOvGvzREf/PfMUFaw/Qrvi9njg8gNZLvrCOx7+bNMUmmE4wduvWBKaR6
GCDrli+ZMHLcqV/NkVBaob2woiDkMqjYmZQVtiV5mQQpR5V/HflNtH6Fu8ypFJbKe+h5WjNvbb2z
7NOWUloVTWqaGOS/197CL2yFm65XxJjvbQE5OkKyxdePKm7z7U+GXfh/7YSa9GgvEpOgzUY5qC3x
GNRLTGsQev1Q0311wiL0So1x2FB1VNpsXddrwHEs2tuPICj+gd7syyOXDUXNlyVdkHEiguLyPEFD
AhfDAzuv6m8Y9FWrxygAMGSpH7BMCl5TwX7VUDdH7ze/Tz05sYJ7lfu4a0DSoRmBh3lC5zCqI/0N
g9/+HBc0fTfsmKcBIr1jieHAm8F/+IvVbhkLdEWqCaT5+Q5nQQWCyxFNzpwuwQsX3bCtDngAIhIG
d+NboNqrp8wgO7OPPDF+ypAhEL0WMUXMNcdnDp6htpUY2FdatdGQqvjoRci1hrYSDGHsv2YXPPXu
8oMT++e6sb6nwIF2zdeMxl2ixkAPfPZWPUdGciHmPbPJM8BJcZXW8QTnbCxqu8/KXy0RiAfKfBRo
MGfMeoeejq8zutm63UnFrzysto3rbrqw2bjFO/YTDuHgjvqVMKWqi6XUjcsTkYlWQPOait8DAlPv
vzqXtlLnDKItolsjxOh+2zcgP8aiXU0BkDkFMK6Lx+Vcm/G87yWKpBwn7SU/HcZJh2u6CQcs0aus
Evj/yiu4BWu0BJFIvKVrRUelkmwYL9tDWF9/zDpoN0twidRARcMKzGpGgLuvkwnEkeLdiLfUn0KG
2N5yDa2d6CaoKiNhDMvH/ToxMzLYRjmmVZZrQrYhJgTH0HQJWL3XkPxVPlFh9V+m5nb/null2a5u
kI2Wc60Dr/Yknp32rrY/SY4SBSONYcnbZGWThPCesSX5u54lSm0GVw9PfSNGw8U3WnLyzV9QwnZS
utyY29mnZ7BOKB4CA4FysU2MLW11oG7ThysewrOADkxVIrhSCtNQq+119UR8+srwOgqO6JdqZhDx
z4SDkp7kEGHjq85g86rZaqwNzAT9inUzDpJ9/PvKsT/2qbUvbVr/FN32ymImZP2BLP25fz/AaIBw
UjgX5NpmyxGKBRwLM6hkmHYEg3XQRXJS4aqKn5gp07CyoX48ZWZoqDbPtCfv2AYSmvn+llz9Nqr0
kx9MzNbfUm5d6EKg+ij6TYopJyb9lGy5P26XgRUy7afyPpXa2aVqflwkHEktLVBl+8+Z2cNA12as
fqT7RQ5Ut24kBGs2ABf1cyaCY2WNsypDjzRRIfYdXRKqcS9mRQxMN2iBBQ1OOTrde8rFfcHgZ2hZ
XB/doUQldbcUof72G3dRb+10cShqepRHgw3jzE6dOZO6GvJZZh2rq7WQvIo0b3+d7jqIsypma22s
b9UWQes52Qs8fpQ5xvLBCGrhCI0j+5TwDNu1/1/Fo5ytlb1tBZz8JZXuonOYoVidLLxl55LtT+jF
CcK+/8eXPsDqro71FrItqN6pxNnS9oRwXqj4hWlswXm4vz5Y0AjzNF+9CcNOGC2lemHdeWlP/MgK
7XDYeFK5T6qm2TXt/Xm++YnO1ZARWQ/5D5/gyytN3G2gYD1BEhyAd4HORiLfms+vnHcHiXYQkLzH
BNeYq444dLmjLk37L0SwbF+OOJIzAy+VNNrwcL5+WWPN2fXAM7YF+P6kobGnOmrbBnawU57rFSx9
uyssntgaf1izwxlWxt31Rv9Tel/7aP6FN2GPqf0k7qKkGATylQX+qt9FNzs2Db+zo+wNgIR+Mavs
0uN6nqqN9zPoRHrm5LhmtaPUoEa3u7m8y4QinXMnFyL7Fw71vRhFi6i/tIGIZxA1mA03Ib3FdHV3
roTEaSGCSm+ivDv/MFwjslGwJdk3vnr4FRwIoYW0pWcItSTG9vh3ZR4K95/kRVb6nv9OfDcyPEe+
FBfnUW2cmjzF+R9aINfSLobeD57WiRdeepbTJ+w4mJEo5KnWN0vFdCt1w78pTmST4Q7HQH3/PmcO
rtMaVoPXjuJQDFxzvaZL2CIbturo2q2+KvA5hMvG6IUT8dakc7hLAH04zGIfx7RzB2snHzFUdLjB
ZVnAiR1ggrX1esi3urntEW8iyGCzWH9YYTMslFT1eaMz/xTwrWHZwwmU/fSMbX2jIEp1PfiK8Xu0
H4/LVOnI7Bn1qunztDW9Kn2VouNASQTFZY4lv3n4Rtd7+SJk/EqdVuG2vj86hEwXvWrt9Ey/+C0C
Nu1PzxTer0T3CkgtId2D/W/zzz3gUP6bXcc/y0o7p5/bEO3hIr5AxmnRIgN0LaHjece/FAE6AtWA
zTtaSHQVgxYFykDo94OXarRGxi0GpB5A9UvAHGyX/m9zcfmcV2gFiD5raDWFAHEx1acD1OGezTPW
E952MU0e47cWaKuE8lBPmTKMXaWF8cRTQS+i+sTzhxFL+noZ8dzzFI4w3uORxp6gxVk97dhGnZT0
7V03Lr+OlX2mq0XUMZ1VIncSscIp4IQEmWGi3hGzWO3m4hqoJ4Zohi5qau6zZX3JH6vDn+mZhKjq
PEthYZ3Jah0r5ALvZpRBo/bVp5iUwYiFvwiis5tYuI1UcLgqmQc7Qzf+piUe/Tr55sLWeCsvnSS0
sqC4hraXIyOZWJ9U1IMX5KZytNoibHH8q1qaR1pdGb/pz0KIX5dsABMSr6P2n6Jh+YvtGiJe/7Ze
rMdTb4mxFxtBqJ73zy1u5GJWxsUJsrwX+ZtG909LFeBXdPgkmKIwNFyprswUc5kZ/1PvVlw6cvPv
CS/B2wZUjeOt/WjkOxh9w+BBpwcuXv6OarB22NAvnY8WPRnzKINn5CCK5uKxucbF3WpTcppT6bw9
7VYr4KJtMB1SMM3oMI8H1QKT+Dkwxky5MSXhldLJAmdpgI3AWWi8x+N7BxKfbVMSsK5/l+0XHVVl
pS9hLWqBge/x17aqlM6GfgRfQTTJoxIhfyVKer/CFjxrGDJ07ZGcTH7aEyJmzpGqBC/9OgHeDjQr
VJP5tSwMmHkHnRfBu0kPd4p2gngJyn63UOiR9Y5y/WwTydpsTYxutThOtKpofP+glueEQfpu3uft
pILYfJ/VRFEyHI70z8kvwB8GoxkFr6V2NZMxjV8LNL/k2g6KGzyFHtgUYj8H94qpn5aIRtkeNZ4Y
IMwr8DfwwK0LzFLRH6UXMsJLeyvNdn6xe2vBHroi1RX70ZEqRcsDeuBW2fXXFkZsztxb2zEXqlvf
HyPfOLJ6YANN1DbV3OkyoII8sZ4zDbAh9rWkcmx4Y19XxWiWRN8+6GcIbI9iFYfTtCzr7Sk8Malm
UNofHHG2TVs5dGxkIx1WRYHU7Xe9QU+xs4ZAm/JPvG6C/WJpKusTexEmfY8quGc/QojlZAJ0gkMd
cUEG8tjNoZxA2ku4xJXcrW9fJWcwOwsdScpowu2ZmLM2dQzPibky1UGd1dSyrcQQNjRUqFao+EUT
Mlf0WLqIntBygJ22qaus1PEUYqIA0DDctKsOX1BSqh8t2Sdkv98qjwQwh1E/yjQbNhrkrTzCeANC
sRZGjDEybdVHfJbGPXakldyxaXZ2tAwGUkqPJw3m+O+gEu4sT9E883vvZA3tfF5b8TG82KN/O9Zf
/IOJet+0RSzKYC7KgsKPJsVYlxQO4EbHdT9noutsZ2g5tnGRP4iUOjz+AQzij8YrG0qhh1RjJcyk
w68EJpfra3vga0KKPVVBTu2Tt+4v/HjGIOHNxQKLpdi/kSaM953BJRQwk3lyJH19m18Qj7/4ye9l
gItk9CaM0ICISP6qQHF98677sMhSkc+1ZjmPqpjZqrEJoaSmr+B+1iIHVG1H0w28cQEWXfIDweR4
48JbGVdjuXyOEqcITLiddpXIRXsS4vtvulLhvqxOUAYs+JnGq//V28+/YOhWDlr/rgDLWhCA5G6C
MqOTfhN6aFvcN6Tsvp0s5FDYladjclbas2ltKyBW+p9EI6wykcxglqnGft+3pNBJoHAki52N6M7Z
5CkFrtcf392nrXwAu4xMkPi2pZGtH4nBWXyon4Y0Wv6XhlaWMsiqILgBKEEQFFxiLli2aqGbmh7q
cQS7o7M4bKBIZBLgsbvjtO6AuCuGoJBUfEP8KbCvmOsjJitx05oP3XjZLRpETTZD+ipU0HqZCD+3
/YAvyv4sJq5T1/O1piqgzOVaMVphh/zWAtRTS1+JXn9g9HWqyRX4fAjbCcJqR532xp7Ta603kXzA
iCz3cJ04U+LJNwXp61ZC468HNdzmTHJgqEW9TVfLgE2n+ufYRUd/4XgAGgEZSWOzYD2f0LtSdi64
oHWHtHRZpFfy/won3weMRvd/Qiwu1WwInSkI5kXrtRHXTUuhgx4qUMfJsgs1OxK+KC8Gbs1w+ATn
dqTFTdVhIfNPfApypq2gEl4UWgas3NokIRP9UPLg6Q1nfKat8YrM4vXWhPvs+isX9cc+F6NHJeBQ
jhRv9xdVwIyjax8T7kvGdoLuF9OQh3QS3OIoyYqc2CUH0G/LeLH7VxYu81/6cONpolw6HB9bY+lR
L5wpX6s7/Zv3qgOKwNNg9r4iUOv83lXxn7BdXe8uoJAgUjmTaGS/kQo9U+6XiB9Z2M9rtlnegC9K
xvbVwZXbO33ocG94DIXSzf8U8K/t55T3/js5EmV1OGesHEYGLV9iXyEKjQiJjVDLolMEabTz6Hco
bjZ+hfY/cOBr/u8OJ8r12UeH5fK75h+qXQq+18oBzj8CUJPXOwBY0rpGvXTn88rAq/jN+kUrTrzT
CuOFaP2KSw/av5KdwXtS0xkdPj+NrEpQDUvyPrubjb8KuetG5HpbWpjKnHWQgou5N/nXgKXcKgp2
yWz60FeqXhNt8unyrbzj0bEtBvUDZwWFBo5E+NZX8zP4nxb9OolDnttmvaR6E9HzE4f396CPMaIY
QddUK+01sUXi2TsT2mwOrTj5nxHLHalKc9SK+xzkc4GOElXWgKNrw9hmktkDWF419s/4LoWN+UGf
fgsedqHKu7LWUi8aYCHQxgx/ZgACqulqD3X23yEtIDLxje1Lj248EOtcxKDdb1E1RcRc/aFtE+rg
J1ZIOFFJkgSVld/ooa+3ij2OXjjl+Lp+8S0O/rQ6g0Vwu1OWpeByGoSUVa/qRE8h+LVjjiWX+8ru
tiYDJ1zeTFJELphuxBbR27i0+VOMlkeiOPSULRWhuzP8cSUSO0T+o32qWfxfthA/Pg0Dp0L69Eb1
hCpzpfUderOpCeXaIKVi3PAjdDd4SlwBJnLPkjKzPJGDEPrvu1iMDP7nUNiQdpDJZWKhYHeGZ3qw
Dz53Rnv8Tr8AYgxPcL1dBtCBvsCDZxrxPspAHjJJ8o562aK3ImIcYenV9O29z3lhD++Cg2r8LN0D
QwuO5p8oQjlQCOt0OPAXyDCxb95KtcLJqVn9PF50bNLBnnX47fybp4p1meR8uS0ujf/qcL05lyJk
tmC3HMo7p+lxaXQ1Sf0Aoh3oEKKdQsvCKtSdVgnszNgHStPVupdskYmkDaLsKJF+huCIpLQQkGIW
upliCJ1g+Lip27KdB2anfArM2zelf3k/IPFRAxM0toAZHUOKJc8iK76KcL7WsMFYsNc4u4MkQN3h
V9GKyCs2dN0ZyB0mMwq+ZkUGAPaNFuHqod/PjfPD7t6JxTBk4iU8sWCqKIfdsbkMitaE8QgTSpxS
JJD1/0doL0LkOSdfkN3iPZfdMBSYIsziKJfqZJ8Tf1X/VtDmbKmKBMVTeefwOPB93vG4MWyGT6+M
Alp6bdSakvq924uVhcpXlCsj2bnSris3/sGlg4vaqW6IZ+NlJMfjgeLDgJWn6W56zgTciMuRyGQE
AfLqgk3ulkjs18qCf06M2UyoSLsV8coabzfmgQFSOOQAjDqPeQk8Np0wENNBBBuJlYSgWrArML3Y
DnldeGmAkELT7Or1NUj87WfKy6s+8vnZgvtkOceIxSOmVh66N8ImNIHTc4kGrMdbRhlq4AtasVYW
8kJPqdkhgBTW7qTpBRxgjcyaRsA/W0iX0W3j5mvY88hm7YUDfZe4Wxdils/48i+30lq18Ow9+2vJ
KnHzxKWSmZBVLsVbYChwBvzmW7r+oJRhCbqydORcXDI0nRFHTCfCoTO6NdqWjCfuHGPbC1Zrr2KC
CROop/SxYwh+/HPG6shrzuMfXyRWx2L7Clji0fPblpgOhMzPSxuLVmTJ3DB5MMfcjptmjesnlxf1
W06KibMUn7Ttl8TVf1jdmtOban0VKVM7jDJoEzTDQSq7XvRsRKhHF5AnWF0akJdilzQW2BXCpg6C
8WMUF+BH+ozinLjcv/iiMpGFfsHcxu0F2y+sSB5lYAuXuraBmOXqOOY9XrOPiY/7sk2R4Do+3SKG
chjv1pLVaseQ8PdcCXy17CvkBJeJxM76SM0vcGZdNl7VA95/PSnv0eyfh1EreqZ6nYOgpoxo5x2O
x0y8CvSpVbtfibLayclNlJgo1toUh1HSwCw5zX4R4wZBq1xfiV73w2Pwkb8fqzMBba73sa3H4vsE
yD7crSS5YS2rR14KCO8dbJNjyLi6h18KOz9FOlKpwrX0cGG/7lQa6E7xGRO2kmuvf+/uU+c8khas
scr3NKnCq+pNeKiWkWGqujdKFg3tX0F3lruldyEMf7OrqfZ5lIpibJ9V3P8Zy5Y7LG17KdaSVwbI
aazrf80ry2956OaJmubtsenfuBVRs68sANPlQIFpwfEpAeT8GiGh6JexpjncHKMpRP8EgCFQPnVI
FNcWgk6JEokOaSk6GGwwbQF/xqKCtPXyWuANJMPjCuoO+gFPYVxTbMp8efL8Dazq2azzHNUGz16M
r9ufsdhcructb2trK5Tgea+1Qx8yJmG6oLFCLIcT43veJyOtlEPte9nLzH6l+oHXaEvMI6vNvz6F
b16dJvirxIKGc9MLhmbjto/ZN2wF38Ilw21KxBvN0Vng7xzgUeCC/7+Rv3B/GBXTpqcOeodNm2T6
ExIUW4SuRg3jcs/TxGAa6rWNb2B57RWPDDlgPrc0S3tmOvm0XWEZI2c1a2cnkR5EMXOsd1PBbVMS
X9E/53XB0ehnpKkHevMeERwx8bKFy0fHG8OeizIGLp2jAmdEHX034emFEkIsF6pNAQw8Mq6QqUbh
VhiOsmXJPlGAk5W6RYLs3rWsbKO+LRLiHYnHTdyhTP3a4R5aDuzpXJRE/XVHPHXL2vVqFwR4thtP
1qBP7HEjRtdmN4xfJeh2mYYNjthyqTlLRSEMfxN7+8caQXhnrJINACu+hnwQ/av8rNf5N20FuGYr
I7ctJHZ0P+o5UccM3GRwQDre98qMPdgLPr+1u+5fASxDTBum6ZT61eY7nVl5GVnkeXLtaRXB4P7Z
w0CI+QzCbWC1GggxbCVfX3AL9GHvuTbyqDxzlnshDrfIrZ5/unfHapUMtdWCx4N5v+NAxJSXNrU8
DdeQqRyb16kUerIDV8HFJBoYZbAhiEJ3zfr/t2vPXWP+1x+NdIGn+ifKLjvgUl0eKCLvsEDf73Mu
s3hmn023L0wGQt4CPPZYMIo2SVTM7R2dzBm0wTEvskRjPfeTAoWNv6QaJ25pp6A3iBTBcLTrlM2Z
JGowozQ3yj8q0n8J5lvUG+z8FQkwZHAQyFO02yXFVWDK5m3e30Jm//aWnd86MPUSAQ+lh29oV1X3
Yv2LDUYzwROoOpV/h7digNueNqYc0HwEMxuC3ICrqyll/3ZLX/Hzanj2oTdfkyYkB9P7tWtRvKg4
x1DmL84ESqY7ieXMWBeM/8ipoCv41BCNU/3Jsu5S3RqfjNF4l+w7R5pZmI3HRLvJGrUcDi/0/n6Y
UgdbA4/PnzJnJN1PlXQwwx/Z/vTA5n9tudEryXtl52B9ZGR0JTOiW7Xr15WiIXYG6yd9pExR+udd
0IsXDBTLK+E0Q4BPpsXAAelwc8Kocy1UuibIVNizRS0/kEIMxo0PRwFARUVhAFeaofyYwxVJodzH
HdJsuSjnL2XIPszNdqj3mqKSIrIHE+akXlceTvmDgBSXEELLiVDrJV+HzxBHZi2H/4d+WVZgBavl
iqWUtHAji1Qni2RBeWPsjPepWc0I3VMzJAqzaEKOb3WisRy0RxATg4LXHw/voX52D2oWtqfsautU
vGzjaFHhp8xWublfJgqr7s70GPnSGwS2Vbv2auAS0w6ier+wmqsccVrD6XLxYETXsoZDFj+Sd7jF
CBRchonXHs7vPNmGGitO0gJY/n09Wd7PnXtqYHuSncZvtm3St7P6CumRbFkvwPrmg8XZsCgfyQxe
jvTey42P1C9Nym4GHb8VsiIrCIwe/lpQsp8+FoPiNVnMtf6Wj7rRcw7yE0aZAaG90gcQbfEfgDGW
whM2l/CKTQF6SOyC9C5HTLrVhL1IrdTBQYdc6PfChfSjDzTOf6ehmBiN0Wl5TWlFA92Wk7MeNWrT
Ci/yJD4kHEVJ/XRe8BM+omTV3a1+LdCX/vQ9PQ6CaSJoejiwx6CgT4f5ZUU8acRr9zKsdZ8f/ttc
F6qdbjBokNt2LNTYd+q6MXGxtNwvKk0Yd7bBQAQbteOXHWaPGUlVEp2/GlgTePHoYGFQjxFhgQ1F
vR3tmr0Ym4ocfbcpfid36Er8xE860Px+A+2pGwkaycNS28SNfCAKVwLMKjB8hU3TYi00VbgqfBnA
dTX9aU6lFXGVgtFWu2NOvqhLqJn0x5t4ppMDcZwUxwDU4cvXvdf0JrL/Y/3UC0SzMmOyMyZaefK4
57m5ajNZuszCAahMlNJ9liq5/yqt/GyuCbzuTD6c3yOXRMOdz7FE27W7Bqn1BE//wLYGyjcx9ji0
B9aee8z86SesKGqmnVp3Iihhq4nVYYMqjkc3Hw1x5glM5+ZMarEV3x34ijpGMfY6Cie749sVwXEd
w3N2H2/tsCvpaWfWNAxmwNQ1cAnuXSjxQrMX9iG+HxdGQPCHS6kwJl5wBU7mVp5xk418r4mumB9r
Bmrq1PNxNuydb6XDaPkhfSVqaMjLfIIn6WsUX4SVtBnJikqsEqQidH6fR3Av0zNx+i+7puceeLAF
WsBb+Pqlb6Q11dnSX4Yrr+xpCm9AsyqdGTBZcRP8N65u6sNsZ9fDgBTR0/OqxzI+rcLFbDQssLUF
bIlmfK1/U92bTbBY5aUHT/x+6a1UZYI0c7RZ7n6zfGWleqy9KI+vq2858/on6voGaJtMWh2Lja9K
XmrXtwAESXVpX3peHEJOekaZe1R/jxeZHBo5kb81bR0dZ8Z0h1z6nyw4D7g2ypTIlWzdSF9nbyLH
3AiAe3/MY8HEGffzNgDH4rw8kdMS93tQT/WxFt5N17zOVtw5DDGrH9FtEED6m9bAptMjbvh2tzJ+
1V8iWsPf57gpuZbk5BEzldZKRwoqep4aPaQVEKz5vFeWVaPLO2jfNa4RFyAzSByBauWUTG4Hm44c
lAX6k2/u/p+7vUyuOgtlWKXkDwExiNO+b+kyBb49ag9SGYdh7KAp4YbO83RXlXmMngmsb5ze62Ik
eZgpFFH1fbaBJrEm6E5E5Cye9nKsRAYOwh9R0zamVyO3xjxvi/Kk7Xcf2ro13IudeRS4vWugQ6d5
3DyEdoe58UqR3P4INl9KmYfDnDYym697kz+xNn9GHlc+fuFagWJ2AkASZ5+qFVoRoQrctislLEEn
qm6HF9qdI8stTnN2HBUKMCVhiOEK1DBLTk6zRGCGjufYRb4Roj1r8FK1EZCLhxC60kzBDoXPFZrb
SA+51gc1lykzYp4Pv+sSOIz/HzUdnotFlOFhsGOxTQdqvnIYh7mUseBaq0RFVXkelbiZvZsmGw0i
+2XlGuZyGD6lno99DXpvl7XIDXGQ4P6Y9Dzi/ck6rHkU2eSN867qJ1lyK/rOeF69RliQqzmCgIth
R6xB3ktBz4R6rolS3O+ikmCoXB0r7sNbQRM+jsG3IWP6d6DzzG+TZ15Pns2LQE5/J9oR52TQ14A9
l4MCe8f/WRs7sjI7yE/GBK/8kNbkvNW1lEjOD7ODx6D7uO51PmZOW50OdKV/vkdqMvWgMDfImMMc
XmkKAE1ifbyUlZ0DxA4brk632hP4DLqrYtMKWHf5E9EqdmX57YPd4bV3jVdtLKSoEBBixfY82mLf
CHmjU1SuCg5qIBYdUQFUY/z5KXlnl1x4iVeX07x6JCTf3CWsRIkltudHWcHatENRjHBe0qqHbewI
qU3cxnbXb2HuOD8SyWLiNsfzkAOpiQSOmv48aOr6sh227r425wEjwxeVG0Sfc4GOZtDfk/pFSSJd
Js89lAITqQT4hQc4IgO4Y3sSiJQC204glWZkfrjxwxPfZ7ZnU+2D29G5HcFlN8lIKn48UVdKuXK3
CJeYVauIb7nu1V1B6/7TH+nN5Ys4AxUDnMfDcXhTLoeVIiXPr3+aZL5yoaCe/+qOYSAiRGfppTe4
/a3dGwqhjeUCnVhfOVJWBIdnfYlSNAsjfeIJPiSniKAXVC3TPEwpARUohSI3lbBxye8sRzpLirYM
cg0TRw2N/5c0/El9F8dpLwm5CEWeTwOHCQFbrWoNRTDnPAgWDUSB8koVQCSREO/QRWE/fh4SHnyL
L5nJcLuqdd+NTBK+oNB8MwEHYIZ8iTFmgXvpgB8c7jMwQRPYeW9kFdrCqY4Iv/EGMzJ+ASGI9JtP
m1YZQDKNmtlXgNy/x6l29g/XI5JfT+K2jXNhaZVFkNXZom4C+X01lQvarvPsn5JqwH+EstpDzkLr
X8amezqURPvfAsu8aiarOrSv7T1VY5ip0nkXTAYu7KVMOmwl2dIR1t17uXSSy1jGsZf3S2+mnMGZ
XVrtTVghWTKJCj/8g/Q1fUDjn1xu+86Vie5qCLAqkwRqNhpl9IJyW8Ovua6G4TU5WeIdNu/ZFnM3
F0JWvfbKHFxxW7bXbw9OI8jskake8wAMvSkRlo807oo3kjejwuzcPTkEqdtcoFSpFxzmg0qKZ2k3
0C2CgFVF69VbZY01gDAsRs2/dnzfHL8Wc6PayvQ2hf75QlNLKjT2R+ShMqPBAF1Ly45G+FcV34w+
kFG85BOrXC1JuyZNq7AFobC6eBM7hQjGrrfnkYhNQaWTwHfDNIX6wzu+rKVtKwoNO8gthSfJ/UXH
IpYy8RptjoHPCoLSs77rzbsFCu3gp53kWSa3tVerSbL0Y1XWObhIWAtqEtIFqwGtZS9HY278vOZ0
cUQkFwhM3AqbdtDOBWROaEICzEBn7vGhwh9EWApVeOVsbpl0M7KBEZIZUwDMdlcXk73k/ptZO/Bt
z7VWRsz6xAQk6hrLCMwikcTNzfshl1pwl1PrIg4ZLIRPV8tHCReMUnqu4bB5P+WKqgOcpuUCAPnc
b5842EqX8YDUQ4sN6TyQ/lWXipXtaE9MPVPJgldSPTYUFwXZityDfZmuP0DE/aMA9u18+ndayFDl
E/p7tQOY0Hfd05dymFamCPU6RTRmeYjVLqkXftKfkNLJ9RR0YVevhdQ7K2oprATYNqjkSEaHFugQ
F/37uiDqrFPwECsssqIdwEbhpE/k2CIbPekmam6izKQntRv61pSywA7fvImteSkfy0SpOGO38IBK
EFvZfSJjL1hpRPOrVlpF9OpO2H/5WGu8unI8b0uWgdh3aZZEXaRMkIuvpmagGK3wCS9OWjt51Eqp
QrIdqWFLnDw2E3OQEznxcsXwMf1OPjJDh82/Qr+9rGPPybF1j/t7+w3LkBiA62KtFxZDxvb20CyC
q6e6+Zz2qmhubpc+G9EPpng8COZlkZNLVZYaBClKvV8oWZvVcgJ3xgRWaV8Dr/pbbwTfZ81tEVyl
qulilUPoTX3MWiFFnnlusOkbz3io1aOC/1Nf9jk0nXC18zF4W4DOE4zlF3o8l5Lmtie1YF/qV03J
WoUhAvWZpDiEdUN+FjHAWsapPhg8Ru8aUmPft0wRbcEZ3jlgve95JQY5DY2/Ejo+AYWEekalRpHN
ye3fh0ax7TshQXqimoH44nRqIyGSCfsGBI6z9JYdOWvYmP3+9rapl0zZ9KR8EOQhbV/Zbw3b6tJ+
1f2JkdmqK/iJJW28FiiVlBsa1hphlMaURDzevDTpgit0OIJJmBxvoYUUygZZTdZk3C/yqzth0aaY
exVJ+QQZdBbFXEePNvV4a4RSNkK70xEEfYN3VlRGs6c/gNsCdLadT/UHmaeTzrd99IW4EH7kbrXN
/X+LFOLhPvhnChylSWNgXus3AYKtv5KGMhbqe+4OyeasxuPQo51CbXufGoyh/SLpId6NmOLeJ0rh
fP2EaS4OKx21WwedGi+UuYKqf9vSzTqOfbROwnkZIeGZmanQyiro/dTZ4pEY7iPM5KLdU5nrrQBP
z/vag5W3aQJR2d4BlrYN0rMGvrbBucfL/gdtx3LXzr2WLXcQpM9atpb/QuRGDRfhqrhffrNPUP7w
nRpkGKWodOJrsDfZSq3tgCoDORcUDsazh104DoKLBsaJoBmh9jFL7rffsdT7CbBmcSp9h+hrLlIf
ZiaCwNhGRZ86oyw0IlBDyGirU8T2hrwfR81ORF2awJhTXh1/oFmNTa5XiZQmQ2XGHHxYNVp7Icgo
ueJqzKQoRjvwQ8ZoQnTpclfP7EhXaCS1D9QXd0esRZCM0SeU/7Gw/Rnhp6AF4AlyAy47XEGLjc9s
arJ1/AbnhKt1uc14ROrnXVoTQtF5EFyTMOT3lrRZSDsD8ePT2EusCIfQK6j7aejwcLs/cfPlaUuN
IFpg+2biJzHcX+7Q1ZTt/bbE+iLZUVQtcTTBXmfZlGo/tB/2Zn10hxR1/R6YVi2KizETjsGagiJd
5xFdJlR9lO+YKpGj1QMSuSbtiKDJL2N1DiYFwalGpSKOQDIIdvMJSI/tki6/Y3Wq3l7bbP9MDXsP
SaZNRV7dok3CAWLOETfuJQ4tqKe+7b3vlA5HMwsQ9RsRujlSx92vSb+gYMCyg10/RlR/HBaE8pqz
MqQ6KQWPkFCLSOzM9hNBqgbqS8fRmTyIaWk74WcfNXNH74XAWCKRT1+EodHPcQoYw5E76Fmpl3fY
yITv9TtcIuxaF7Rh0o8isQR3cMwo8EINA911Ay+/f4jDiSJVykLgBduz9X5fsdf1anfwDpW35BgO
Scq4JmNvAxW4iah5VyMPyWHd5l1dG1KpSlIQ2OMGufA45HrRnq9bQvWR78QniLa+WH0gPv4GGcSD
KvhH8/vf2Xw7dx5FOCcN1XpU6SHIdfIgv2Ktzdc40SyFC/XXSOMm978uidqVquGoK/U07aEs+RVB
e6PjhLZnVdY9i/NySJmBSqoURFsL9Hm8YHKa9mXWtb1xP4f9MVJshk8VC0gcAFnUo70Bnh+OP9Un
cmYsI8VfbETpX5zjPcJp6bYLCvVb1OQHuay/0pNnzg7GgLroid4BShg1EcXW+yQVlf0c5ZsFivdu
vnBITPjHUa/K43wh2cfSfQB838NmSpJsTD5twa5PS0wXsWlmeaDLueG/fCQECN4RBLwDfMl464+1
8GnVjQ6VN0jDUXnb/j3Cz2N81bwWWc+euZSrLyk+Dl0huVfoYy0fleih3Jkt5Gj0yXSwE9J4NsC+
unb0b5+RzEMDPCCNXsINi7oTBR57vAJQXkLOq2B44AZrhk3QQBAr0FMIKXVFBrJ+cjhwjEMzm+2v
wMGM8Owo11EoX+CDz1r8tAulI5aZOQPXyTOtWzsc1e2CmmSiGnwnfzv/vby6+ZgKup5cR+FAiZ//
54saJCHVWK9K4WrpXDQ58sk6KzMfjwSnOAp/eVARFi9tN+rjEizeD1KWSyUaToeFjzs8GM/vEmtG
7blZSWwdfS8ZQH48r/P7IkrioNX91aw3SnjBQruL4mjD6b9XSaGJKL8A/po5SOoXiAVcGjj/5pTp
UVVzxxbXS8XddsJKTom/BgR5YWvAaFHHSyZK4bGYhK/kW5e7Jjv8HMcAHCRXyYIrl0IZviCVvUfo
L6qYNSWYExhl53xSif+2tbkUieG2PzydVb88du3DtkQgCthiE1LFeONWCASpiCwPE0By27dhKxPN
CkiCHejni4SiTWOKl2MfJCgcUE1Hv4hPyeFYRdJ+bBOLLV7HrFJdJHVWQJwNYjSDmrc33237mFfj
9BKQzRYWYVIUoGFE8Tm8MkGeZuuBWCe3KTm2FurA/BxpV89fq57yURySqmQjHGe6YZHxp2H7JtTB
d6ks6gvYta9v2CMdG80028iZp0SE3N0+w8NebE3xHj3+ztK3RxJ44a3LOwkTUTwgD8BI3HUfvdS3
A84y5KwJJI/Mw9y5zfxmdGQl6GNOJp+ATkjRz4+D6H1UskbrKjuIINnwlr665DhMXxPobAL/tMW1
R/PMrr4ZxxgfYGyrjU47crwHGaJDns/FOLYL5WrJ1HuyNkYvoqM1Vl9l3emvuQqkUHYWWLTOxSnA
JXFSnjEqcFte+NDdcPiEeVPNRxuHZUKZMa0eqC1uBgUXhpGEA7myckr8Eyw97s29IiDihKA+rODc
V6qnJsL1bh/gi+PLbps/7+5Mevb3sjdFzJdhOf2pYWEeYaapH+3FmMpLVL8Y+cQ8wFDhOsRf/2WG
gxY3kXGNOQdM9vUVgOpZKiVFpVAEeA1obUfMq1o8WzHrDVikYGo1uqYzd85CYL18AVdnb4YjKhGh
6bV/y16tcrVtho1wD0NNNEiP+4ArwpyfWnsVu39lhzitNGYfKq3NeOTr65gXJlzPnAj9w5RchMoL
rSXMcuJzQGCeIxwESxvuaL6SZcZXEsX+ArFqmzWMKg9i8zrGVIApLwRdy8Hh32/f+EbHZ00m6+en
aNUwc6aNgoOKPHPJiTv48PmLl9MbWIwvF4I2IbV6+U9F4/yrumQG+onRklge7fd52mOwOQm/sp8b
rp1IOT2uSu7czDpj4NRtaCXaB0HzlygESm1jsyWwfofdYPn4+vAahwGQOLGVdb3aPskANJ6kldw3
hu9PdWtmn3ZGquFf7ax2bITWiYb4v16QazUYiBHuJSSmEHjRAobwi2CtCFYg3LTM4OzHzhT93Iu9
nnseprI9U4qczXupb0CKSwnZq6ybMJXJiw1yGiPFABrHsLKTmYOItk4n9tOxO6X59GXCIlC0GUVI
B+uCIaTJ9V06Ozu19KYe2FtzImlI4gLdN6fd+s8nSLiLUeFdhfJPOhkkZF6/O+FozltHXYjotTgU
8K55VIUzRPLW5ptwQAS2COlxRp8nTWjJ6JbYdPEfb+xpqEq20eshmLqI+pnxjYpN14JmjR/0Qa1U
so8Wo7qw4Rmh7YPQnEyvzmVUVmIQp8ehuUdjlXpRZN+q/ECG1YAlKZgaWWBhxGWNvF45OmvckBnc
5yF7At6INaG7MaEkhT9t3KK0BtLnAuGGiReZ/dVz0/TNBWlN38xJc/u2Y0BBq42yLWbnn9y/fulQ
ifh5DecKj+ch4uteNRPjObItNs+4X3/EqdFpAxwI7/T8VPgANYzeCX1wtys13JtJwMnzoC40Ncyc
fWTOaS+e1+dw0Z12SWVZzfI+g+X22ctm8pJNQnby7oqvGn9pNh0r+Q+WFRiE4Q9KKzAWPnmMRRWr
luMTCgsX+vCzyCSieYRxerUv8r6t9S67EeE2EIjit4hSKtvdaUFmYuJHz7k5Se4ILpF2K/xnuhbn
lSjmMhWguJ12rBGZE05Vj/+t098wmNoWWrkgY0jC1PjZ5sJ35MR2fwWFGDAzrGBkcdgGPX7iNso2
DxRc3C/OsRbxtb+wtdIB9pxtgfYWpg9UMy4jcWTJAvRWx7d1u20nhqTDINHk8DLXEA5N/sApH9d4
EmV5+CwDlO1DHZ6ydsTFcKKhXHOJghUu/0OPfJQINiAouLB49rHFagPtWk6s6Kgu7A8e9N3HaAuC
2sVOO5T/rVOcGS4YlU6Yq+ERHDpRIL62avfkJZWgOpwuCLBO6Z57HXHylF4B47tmjW3OdOysbzoj
HTofEg+oyfBOc+Cks8DA6IgOBC2jmd8TN73Bkg133Gipu9uJR9vodGSfkqyPeRl38E6yZwCAptlA
VpKWTvQ9pkOii7ajh3J4jk6b+FD+rj3HTEOwUx/8rDIQzJUQ3LfN40ieLWbZPbOXD96OZxlbkioS
NaocBIj5CCsQ9OXCmrG7AC/AJ/8FB8yzkuDP3zZhjFrqfPfBb5O7uD+gvDFfHUr0ZsOmLBhqYvIR
uid/ewoU2+LHMNsVbT1xdbLNdraFCdBAYj9zHn5XMgy500aLH3HaIbge4CUWlsYcFucmEGTwricY
RnRCpYSvpimmfuXn7UoGv1/275PZCnAZEXgVv9Ef9kOOank1hVHeNWC5/oCI32Ju2V7JjcU8+Hqj
6I7ILQdLt2fw5Es0oaXGWvCWRhg5OuXEB8iS5lVHHw5NX/MHHF/CVC2bUH4NgmLbf2Y8BsNRxx3K
PzK9eKawqPVA40YnIkNvJKnyBGUJ7/GWO2zFe0vUxvaRpyKQEkkWnOqL3HfhbiQwjDQI/LB749dI
HWdXT7XjLqYUdkEoblAFaurADRkc4aWnRFwjGzDhROT6V2YNIaGGHPYgXVfifA2AAnKQfmfQ/lcU
0eLRuR7aaalGZfI53ZHz+C1c9s8iIAMLzh4GAJ8f0+wx0xvdbQiMieQNcG8hEn5ItX+T2hkxC15z
tRZ9nCyZ829flF9qHrudL6uInr7WtMpG+bKiRkBfGgbt5lEDFDDqhK7fYBjLlpDf8wd0KPg392k2
WMicW0u8AAmU1eCLeaMqsYwBIGviarYj/JjcqJMZEmnl+Eh7LIFnp2pXXis/oDlQi2s2tx7fV1XP
dLYfiYBpAlW4u1gYLPG7Pq+7dcNi9INxrdSGC/4tcTUto4uks4vw8tDgwYa8D2OLqXUmJsyYTpA3
U7/Fw/vj89ZSw5o3ywALUbtjnOC9QowSYG04AfWy1b5Jv0rp3/itgm5auTQyvklcJ9Feanye1Fny
9YGT73QhprErc6Ccax/VeYTsS33YdbNbU1nzVMfEYWdExEtGzCd3QcfFLj8Usyk9pAP6uClkKI5i
eyLDuVAAcNWAuL4p2+AOplDrb3IYZ8fWNNJSw08Scj5uJtD+sBfgBFxKtfIWrQw3n188UzyNQRet
I6NhO6E5GqOrrmghWI65JYnkwNVrH1jfhJ+rmqvk6e9H1YA9cGApuoHTS0AWUF1IT1/zDYDS0xOH
X4i6rzv7Vy0QsjNnPnOeBvakPZu1It1WZdRZAuuvu6oa4WA0+8Y2Ng33Hp8jyII29++jtM1LdBaf
dMolZt62EhVOyYu6D3tZGI4bidrEYQ1QpfmMMe+00FmgciMFbwAgXRt5NoXt62WJiPzWpmfdcv96
fRM1pK0BB0L36UVhTfmw7IR8/0XR7Q/LXKmCUrWoHXbQT/k6A6n4hlc/LIkFr9iPO6kfDgP+zowu
UOcObKYLVM0x/CFn/2M5o5mFa9baTjlIrKgQNP8tvo0Ue1ApC3C/GgVNpXTWhm8QVs6v+H7TuZVC
9ZkvODrdbUFm2IrbSxXQXhVtD+NXbBPzwfAnUvsiZpSWX4Ho988wQ8usuk1yJQ/ZldQLKp66VUgy
jQIJ/WU35SFl1+T4HB69ZO2tp8sbuROO3lUPLKd/h2dct/mbzPjVqDg6YrvRXdh2WTdjXLL480ch
KU9aSnBnJVJ/xQ0mhZjTzjN24xyybnN4VYkLxTm0WT1LgWD9IHGQbnyrTQW5Vw1Gb5lKWVdTilSH
ReiX7Xlkdjci9nRFX4aPLci08uigD+7w0it/rbK5sdt1e279o5KAIcQ6i9m4Yqnye4pQiqAunypU
4azBxFzSdo4+bGJpoep6RCSZIKk1yfspU31yj13Q1OEmdi7X55kh5v1QzgFRFnWADk1e1+NG2Ekp
clveS5NOKhye626w4rX4fFclj31YwLAMfiUE9/jYoJcj4uiFR+ZVHxGWY2BYqdIE+iCpLHeScmnt
bZCyK9/w1duI67VR/Ytv11doR5I1gADVQEmAVPw89+tXWVQvbkBmEmC/ITOLfONFiJQmHnYUUzp2
Fr+8moPrx+7UDK+Bm5JZKzQNGm1pyfNfH+GQYPIjc6XWChaH6tYrl3V1IIsEvIYXl7ueAwIAmDbl
6y2s8ZrQ9oCC+wxlwfkBZX0pbmzp42Qh/PwsnGbvu4BYtVa7tQcApwfAC9Ry84O/T/h+XzyVjoUt
sYnxpGMj2P6cp19g4aDq0jnZlZ+imOFw0zOVFhg7rcVkaqTU1l2CBO61kmGfi9quDymIW71KPjPC
7wowWxcMCft3ZhWLdD8ipB6oP79KaOM5zhOlx4aUFZykkIqF3RSln1AYEX6VbPiLQMZVBNYDL3Q5
BhueIXFbrOkogeueGA2ZQYPj17awlpKfhfJ+x2FnKnFRMqWO9J7uk4qo04Ys5NQfCR+w/z7oGh41
y7MUD0E9+u3nm9cqb9XVKkBAMtFLTEIjJFsBth7sS0lA1mnGyQ2zSXI8dR4KrbNutKqlJtT5wbbc
DEccvNHR8EzeAt2dLDxnecrJKJhHcyzBE4Dry7u67gT+L4qjlr+sKQk6EcUjaV4npKpKnvdNwjVs
1vPCltwrmbOpFKYao3NV5+oFxonj+7SrwCRW/AqGVj5EoedoLI4IbF2/xSGV7qS2QzmvhkA0om9s
z4lBqktBfJ5wI20w4eOXUBpWFHf1MAJIu53ReNuffDg4B4jwkq18svQAerFqMMOTO0QBjfX9MYJ7
/kWrSyvQJESAGpHAL04r4NZyVNdR0AOIQvv3tcq1nhj46CQ89ejZyEzwveubAjZk3b/ihxDfAdwX
CCkW3aumvDHhYpwj5HyAdP39RAl1sFwpLkaUINjcVTjFXTYGySygmhpVBGiN+P4eRXIJdBcCAqAI
1cp4UPC8fJrq6Vdd5n/wEzVIoFdsUCGM/EmLyJgOyQgjyKt1zSFD9rg6nRUUudIEuuIhwdc+QnkQ
o8n4h6YAi4YbUbOXpOJ/mOQHwN4hmwHN2xgjYGCADEDzkp4gswvPqqzQ+CBNwWNVq2Cmorzqffp9
gU6P9L/VwkvJnxagMCUsVKIkv/8Idtd6beqbGRzS+7xMc1qRkI9X/onc7FmP8fe1velzjb9yVjQp
7pd+/LSpczgUAGfqxOFHfrBcAxf/5rmETYm+MspWxx2LML0N26jjpHCQrwWPyG1O9B85TlJ7GCiH
yqp/qgve/PUcY3uQLcO7u465Y/F+yj9oxtm50tEQ4Q4l1SQKamsH0E6D1zsvRjLhJIvqLhSCjI6n
rBfdY0HYDfz3kKyNmtGTp9+G0mv9PS3Lhz/platud30hPSAkLkDNhCYx5WtqIbb7I4Jh7ODge3qz
Dj80+yMmK/82MHIVoHxmC21zoYKfVPaYjB0OdMtKh5XFsGfEhRm+EV9qgZz9AneXzsQzTKBC1IcS
b9yqjqo/aFgZ58GUtWI2oVC/VnRi/cec/6CUJsNGWMfuo6Y3YT9uJ1JtjBOxpDWy2G8Kmbasup78
bHIZ5TNvUj8p6RaZhHOx5KF560Ey78iOIBAKq8XCEHqVVSfw0Y6EqBf/I9lS+Bux0Rj7evmcM/wh
cnUdbsrBXYWa6z4VX0Pp4xY4auSeh2sTVq2AGcUhgKCt7jwtB6N+N/C1WLU0BCUeOdi8j8aoLjc9
s6kXaEi8ZYPZqYkyveeNkKg0R0q0VVLBH9MHPBpxqvmxDX5yUnMnj5s+XYGlF3dpkqmCDF891e9g
oMRW+21m2nbD4R/6ozhwWE9Xdx93t+IPpuXeu4jrLpmuf4BTrgXFGaLJvylyu+cr21Q3X6YupMFr
cvUDUwUuqS0N2TmRa3i3NekbpMmS2Q2IYYGfpJvC2Noc/RuARe61DZP+O/sV52G/nFVh1cDoW5uX
6Fbo4FqmT0WEPkKK3GbPhzIDP0kqmnE9xOkYWDXSC/lkWZc2izgRQNzYjRUIsKPcW1UpJo0Bn2PB
LMRNTcYX3/ouYBX5p2FooPCQw3NRAHUeev2/lPSTKGWBVikDXU4hPFKhi/bHFxGJXp9kbPViSjka
Ncwu5oRxJOBqCZREwB9eYtDSVxK3jbJVblw8op5LbvOzLC7+KNDGhawHQQc3JlP1N5ohQV+GvUbL
s7FPNbGRnfV/zY9jnLp+rY0kG+S/4QhXqqQgA2ty4ILNr+ij3wiO2ApZsG760OtlJ+FOMz1ZQ0F6
wbJiUyrVW3mIk/ti4xV4lC8ZhB5mqclOQawijlxia8OSaoHAsUMUtR5sS1RhWCgOCFuVp7Vu/5EE
vxQpnvkjYtYhhO1+xQBHYQ1NX2kpkxi3u3y0FDDsUFsMiPdTlJ76ZY9WoerItRNVyeN0VMF95ArM
cmbXGIt+del4H1OpAAfZNy/SRQ9CTAxAHDNedzHOq5LInRdpcSlZDiuViY6Mo4kMWdEQKoXVYGgL
kH3tY2T7QkQjylZLGhkjujuPahqu4wltbDgZxa0TnvffwNjFi7BKlSbvLKA/zqZNZbt7z3ogTF+M
4FwonoO8UHq68Tmjej2rGyUg4R9JTcrIy1zJB+2Bvab2Yxw8pTEZ89RhppWgut9hYgswW48S1IAO
OZtRixfjMSXZ8nI1cwQJQLQcvofdCcPAezxas3cfCBpsC+Y8gtgoWVKvbT3lwC6SbWHn0oxAFr2W
t972KoGPA0uY7Yh0SthUKqURO9DHNMda1nDahu2CY3TPewAhJBgpxHknqIV8jqy8zqDQ5/5z/KVr
wIpB34etbp+UZl2JU2nmi28Eh/JRtQccJ0TpIVVaAPcPtTP+bVud7x2sd2ab6urB+BO/9OPFblP8
RSeR+mlI47DuzABRFIIBIFfKjEX8w0SxVqx0OmUaKKfmYyjwrnJlhq1EaMFLqML3H10jX8IJUeLU
uY8wlVEGxLiisxj117YLMKvaUh/8IyKTe4ldS7A4bH1C9nGwF/TpATjrfJJAP+3HoE/axgj+Zg9Q
eaylT4miGHNsgvtP1PgnQHtT9bpM+LBVLuTOBvQ1hJoJaSAfmfJiq+PtQC/orCcoW3FxRB+PW4kR
esUbGX8OIrtJXbuhbHXxQpLOtrQMsFT3r7WO/ztanv8zCtfEVyf6vCWwD7ouC721sAGxbwoKse9T
cCMcxGGB2O0nIIsZoSsHSPAjn5SEEsTrcHfNdRRIK88+YH3BNCv+RBoROQ75GEFHoJQKCuxW0pPL
1wJg8uKyxVrHQhn6DA634CUAjQY6nNZ6rfmG2vM/r7DZfn97IsMUk+Kw3CSrdXxZQ7o7mAw+/ADi
+9ecaTGocJpwrhz90JR/5XyzwwXEhmFN42xVauX9XVMO6bw0coOsonK1UnFmzbxatodre4JZxmSM
S9a6+i4loae8lJUFwA0+5fA1zCrZen4Hh2/FZGuZ9BD4Mx6OcHsMUQ1KBLUzgT0+VhIIw3NAIt4l
GOzwnSj2ZWi+hnPnlp2lwXc4y67OLuwAxfKflK+JuAQtzSyjrdjxREZ5L9CWm0tbEf6aXD/MKSTk
YOpcVWmmv24m+PtLzfAProSAj1G/wvOjMFbxDbbrchp9Yjs86rqMY2Tli1OkWPM5UYB/Jk/q+W4N
jRkntoexhqJXrz4IamWdTBu1P6vQy0eJNX+IRcgCXmoqmzBu2dMN57tVWDJXzAvKfAODouNkMPsa
sJN+MSfxiDbsTDNVAhx3NORy+Gku90+B8rZQW4+/BdOlCdayQb39BJix2dDRf5OHI2yOhM1iO3Z9
fk+ZrN6GqFI+Y/dNgRvDjsjQZQ/1XPwdzKw9+BaRAUsLdzOqvS6c5WjcSbMJZjbe25RkMGwGMs4h
9DOEb7o9T+u2J1E9zc+zRkAxzYy1t7XgOf+E3OxhzYhmJ0aV02nwREYypNCE99Z9QoKdSjshVcPf
BGkzdIH9AXSKnKbMcqFIHAVOeEWYPdO1OSV6juFTgTK05FOXmIj6KdWOagSzgqA69QyIbHw6KKTs
7JRENabfVpEEClHQSjCg2xqQCuYU+7nP8SNuhSr8H8K/cFS+CMH3syvXxn/zPBbBFnhFE5wJPecI
laW5sFPl2nbZWajmAYziIndlzH1VzFA90Xk5x3HPqdL0DqzhyEVVjpLzxl+iCYK/zvU7EGo7s+Vd
E6rp/KM2O+04ZNMo2Z842DLGFlKq+7RKK7hhZgboVRmBe1eJedgkIFID3DO9egI0PdS3byQlkT/D
0Y69Qj6VouLdvKV479q7RI/NFcKtDQLbC+BuQfADMWN9cMskJqQ929c1KCIuPxu8f2HHfu4uGA2B
koHUm2HfB84E1hK5byaPz3ovCFP5L/Qy6uUZR5/3DFa5mbgzVZ4z+Rb7zerATs/dNAWE5nyTs54c
kSbNZAcxczaPJIudQdV5p+9KasMqF4Aw84SO+sYKlVejF1Ws4zGq4Y+77QQ9yZviKgAAvNK1SaNK
kb9wfw1/5l4WXzhCm9SvI/IOjHkkAwphgnaDlX1s6QbK+4+qBzn+nRsHg7+yUzMCP6cQWATUulEw
a6Yz8qfuUWMZrOZ+XiQNVyN2oU7RfBimPnjniKLY2YRxfbgOPNe5dTX8Fh89DpdOQjWqSxe7f1BZ
qg+PQO083I7Fu5i8MCLnRPqT4ApBMNelva2yD5kIZVLIPzGF6JvKkuUzVlK/hiqj/+bqjaOU4uU1
Nphtw4sYWt2sqkdgpQhsThUqfhVFdRG/gZWQwh5+xNVU0g32pTrJJTEmSwx+khYIFC89pfNJxxE3
Clz/6KONvfNm27RB3jti/Qv31/dz87r/8aEgNqMsev2WqR48qtXOhbpTNd/Y4S5jwu0D4u6qGf6B
dAtX/gRhxIOamsMTxoNSf5t+AfceXk9WViVfxlD3BQ6cPYra//oK5CRi500KyXtT/9e3ZyY8GrGP
HVLgt/A5mpv+yxu2kTepSeEeVB2kvnfF/2AW75s7Pn22h7SW0jgkppVrCQKbeyqWW8XeSCC112Aa
OP/upCOFREUZ8hnSuJF+U9Ey4T2fPHHj1Vr88tgcouOdWQNKuaKA/wDetwcnsUNyAuan8kHmjE9x
u8o/L2k/cMO0HfKG2oAduEo1Z/54GmCSDSMdcP7pm+/+gmigFge/5cu6mcka128BImB0gD7CPPxa
S6K7N9n/9GmMnlM4z/NnFBPq+OQTceVxBGE33fHu8kEaISqnO8pbumaqS6DMIpDXF3sj6k40BLLJ
v74Swq1ODk6Jnv4XxWl9rNT+HEAsYqxgscoTO0OCy/OwQfYvOHQ5BEm2O/vgkDbTa9ORjhhuJ2Zm
/IwUN05WvrnCIu/AjEn5WKhN+oV8/LuBWEW28TkZOq6hv8lvCE5sweLG9g/hx9kyTV5iLpIxTA==
`protect end_protected
