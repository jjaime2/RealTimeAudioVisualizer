��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊\���$�?�#ظ��&H�%�慩T&�w\{)�eΊ
&/����$k�p�z�E�0ibMe��3"����9uP���U���;tr�VDZ���1I7��&*�/�<I�p�qn�B��Բ!X���<�<��
|�}�m�A��l���+�o����]#R�� �EHUN���9%��I+���-G��ii"m&{�O�`n�iB� q7��`�̜�R��>
<�t���"4b���'�QVr�״#�9��u�_&���g�!�)Pg��W��#30w��q)>"C�����|���Dp����3Vx(?�ַ�)�\�r�PA�Ex�A�-\���"��������(��DD-ʺ��f����&�2O8�2n���n�h�粤~J+y�	%����ۭ%���{z*z0�����˂Z�u/����\��y��3��u
B����E�q���i?���'�Z�'/,IM�n��,��s�� =Ay=�,aG�M��Ō-J�3�[������(�!�D2_w[��5��W�C��O�����I�0�	âte�U�4i�o�/G�P���#���F=vĜ���q=CC~� �h�Z}\�@��^����W+�m�tK������3n�ׅ��Λ��J�_�J/Ʒ}����!;����78��Jaǉg�9P�Rcw+./�J,-�z�6~8��M�yI��g�"�Pb�)&*5��cvN^Z�3`�)��&z��xׄ����8��ߊ֚�9睴K?�ظ!F%��"���$�s��zE��'~B���;8���U4�p��S��t�Tg�es��|:k���yC���LX�6�ґ���֭��y8*#^�w���ۮ�b�5�����t���R��G�X�Z�=�@�X���|0���YF��{>JX����f� e'v����(���+L�/*c`g��H��@Ӣ�v���(��15s�����m
�1A��ް/h�ps+BK2ƫ��\�y��gm%�T/+d�l�i������$���+���H(��0��t�*��*�E��A�	$�t�:]�g���F�D��%��bLmܻ+�a��P� s@�%~�.;P.���p�7�?�l}�8�0w4���5W�	��L�M�!S**وt���<����}gF ���}x<���/�/�є�Ic�����P7�܏9�0Q�\HhS��f��L	���(l�����s2�ʬ��q%"��~&����l��)
`���W{����uj�UL�C�?J�7�sдֲ�����H�)�~�+�<h������:���'Mȭ�/ӂShBa�!��P�.���b�m�}�F������l	7�؆��ֹY� ��\�(�]zGP�R�3dg�����e{��K� ƗChx�����R;?��Y�����p�@��L�����Qi�+#q��_ͪ�	�E&���j[����]!��8�����u{(�O!�c<�:�X������i�hȣ�Fk�K[_:ɐ��u����P�<���m{>6�;���G���k�싫PM�pa[�a3� ���{P�j�6%Y�}}��C�f����8/�G�{���jp�I�/I=�"��VG���/ThY���jG��8�x�٢9竢s�h���9��7�;�Z��,����+� �o�T��L��o�hEzu�,��z�QPnmU��:�d��$�aޑ�~4��%b�T��-E�(	U������O~R��"�b�s
K�u��(��9��]���Җ�<����.�d@}��/�b{�	"�A�Q�'{�? �As�1��d�梺o�0p�ñ�Q�MW�rR��ϑ0����c�ԛ�%��N��Ϡ��ŹHbA��ᡆKr�i_V,�μW{7�ӻ״��p��5�.�=N/�g>��3F7����~mey}>�}��(D��6Bfg�� ����/���@}�u7Ƽ���Ag�@��#��j��6�`h�{>�2�9%'��3��f���j1�p��GTu�S�j:�R���R�J��Έ\�g�H�.�yؒ�29���0O2C�e�[m�=�#Ib��U�	���Y�����R�盌1gH��ش��!Z�Gb��I����wۻ�X���s��ȸ	�����U܀��`vs�Z�����B�V�Z��漣��� �z��`m
O��	!-�F�!�sd�ϱ@�gJB��[c���I�w�6<�P�G����MWQ�7ҬX��o$.�A~��++݅0)�X`���A��S�.�}O���8�.)^%�gI��j-u���U��[X�2�eb#�\5�#���ƛJ��f~�/�v����%���%�5�,}�L���57�5��x�z��:���jA?�C��f�M[ �(��&7�7������w)�Ғ�����]Qq��C�e+e�1V\�*6�FHp�.s%(A��^]8��31���N'��wEĩ��Dʆ,l��'oō�`��ƞeՃ�2##���S��,a���<��E�49�^O�a-l�^z"/lt�"�XT̸: t�@�H*��Q>���_��p�YD�{�ʗ������;ПJ쨫�z�痉����'������W����>,�C�[K��W�<�<d����u���@j�*s�L҄.�aR�5�&�����x]FйM.)RӏGf`B2\�w f3K�Hz����&�$Tu�z��v�Ġyzj?��ZĘ��`�v��'�Π<^�I,��6�yx�����1(������\��+ա[�b�1�.��+s�qBp
9�z�=���} Cٿpr=�H��~JӱP��@+gs��lv��a�]+p�L,FKoD�� 8�q5�ɩOt%
j���&$+e��'�úrdd���3���.�]���������IWջ��XQ��阅ʞ���4��%�������/$��`���b�@��"��xt¼Q��4V� �|���.�W0K�7�z|���/1��'�����9f2����p�p�nx&nL��H�4�߳]ٔ?�u��}�u��u�ݨ}_�������.�0m�[T�<��߭�6�?nړ��%B��ҕ"z ��\����ob���	"9*XP-��9�I��B�:�~�%;���%�|Q���D6A�rV2Epu8C�ˤ��\ѯ�?Z��}�o�������g�=1&��L|�bO~�	���RT��K�/��-NI/a�YSl��r�-:��V��2|d�@��5���������7{��{줹H_L��D܌x������ ��xҩ�:L�x孪g#t@,���W>�ě�PV�����yv�����~�n��Y� �=Ĕ6
6�6_x�p�z��5�`ڹ�a�pl��D�d��f(e2)����hE���Hk,����J�41Mf��� Z�E�Q
�KՔ��$>>���w����x�P���Ai����mW�ag &"#�����c>r�mЙ�d�6j^�rmP �F���ƕļ��5��5g�p,,�!l�%��+���ח>%���Ѯj��cܓ�NƟ�w)���E��"�\ͮc��: ���"��2�O���)���#Ct��5��rd��9o=�q��(Z�	n������@�ڽd3�� ��ڮ�X[ z�z	=m�1A2RM����7&^F)���	���<&Y��Й+�Qln��MA�6����)�ъ&��Oц���#n�΂w�d�cL�^գK�����19ׂ������Jԧ�cy_�.�)�,l������킁��G��n-�x,�G��y�����3�<m�P*)&YN����Y3�L����o�,��� i����;��+��1��������#�L�$��//Ň�K@H��C�a�bOŒ^D���W���{>]�_��� э\t�Re����4BPosr k�4��y�}�%'!�^��G6��m�!��9�J�8tïj�TUX- �,������v���Q�[9��k�3��Ĩ�9��*%C7�$��̿��%H�֐Q��N�A�!4��Qq���C�!ۑ�:S��p+B�M��B�Z�#]�O���C%�AD���9AmId7����X/�gxO1��&!㠲d4��4�;�s�v�b�C�Ĵ�����W=#�/�]�HÝ�c�t�&�n� gF��"���j�-�YSTP����6��{�8�iE 03�qϗ<Y�Q�n'�y��'*:jJj�*�гn/7���q�T�C�0��\쾔|}����`���H�_��Fh�C�m^������  u4����'��ݲ��vܠ��)�;���Rs�#��Y������ң}
ir��
P.0ף'#K+�0�FNV�[��XbGj��l!�&�u�,�P%��Ou��\�;�w��a�qp��p��,����&�����6\����/eG���Ύ7�^��į��_���S?�v�B]�ۍ78��x�A�����-��mv��W���ȞR[%ո��`� Aq��