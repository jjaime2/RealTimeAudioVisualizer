��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���B���Э [$�V|�|��?d[Ѭ�(��7 ;�gG�����h�y(�I��Y\)VYy����Twr�#���e:o;�K7s���b`.���ݙ�%[S&eb�pJ�J/a�Z��W���M�s��&��Γ`:��57��9w}l��Hcؔ�T���M�z�\B���qXb}-�m�E2��W?�.r�0"==�v�%� J���%}@Q�\������Q!��:(�P>��c]�22-}Ъ�������6�m�Ґ`����vb	���׿c0E;{yL�]^�S	�3X�H��=�<�C+��C�M�K���OP���!���űáJ��C�Ź�?��)���r�,俚u<�f �R��-4E�Q佞1���:�]�_9�0��򑔇�?W���v���N� I0Ǡ�j�ƕ��	�n�
�4!�d��u��D#�|��BY�eQc�Wk�Z6�d���6�#�iGƏ�_�s�9!^�h��v^��.炛0w�2Ƭ��Wp`G�]��	�{���J;���wA�\O{������VN�{���@8����p�7��]�Dt{�]$��l<�������0��\t�`�?�9�{�z��_�VZ�R_�.I9���\B�$�t�.��IO�6w�7�㓹rmv��b����z��U5Q�!�\,R��9:�o�3�ګ~�:
ɭ�`�t>o���2����BI�w`8�~��r��ٟ���d�:b �;���|AI�\-��-7�9�L���vF���ʻ���^�<ܹ~zH���j�#�����X����qV@A.�vj����A7#���ǰ�\nn�1MfH6�z�9)�ӯahqQ���lퟁ�'��f��7��A��2� �>�?���"W>���@�dc�E)�,|���Rl�z3�����ZY�C�^S.��)�}�S�hµT�T}\�5�.,���)���$:�&�)R��?�(��,Y dh*+��KdN����=C����U������S�86Y
��E������+�^�T=,3���$aVX��[��1E(�W|^i�� "I�1V�c�=Ĝ�W��o9��&o�³�������UaXfS����d��*m��]<<x-��(�ʻ�ۄ����]��bԲ�d�Ŭ���%��ȴ:�J?T�_���y�6~���E�/dσ�����(���mؚ���B��I��3_��;^ R	��&X�o|8u#8`�cHs�ְx��q�ۆ�r�|:�Y)g�w�����Y���fm����`<�P��!f�>�����%O���`�lvgB��?�E ����8��q;�[]�7Ň�>�0*��x�˪f�T��h(AJQxס�,�#$)�]���H�H�a���B���,�3���?���iA�[+R�r��z�k�7�WS��wU�:��G5�K �|�.빐tL�ZU�sʷ-:UݯG*�)�Uw�*:ENb~R��3d�ϥH�n���-ʨ2 N1�HB�~*Q�l
�gp;��xV)C�i�KACܓ*����]�h�@{uꨞ����7���gMd���=3�5���{����g�\B;�&���k� #Y�������ڳ
�H� �1� /(�B�k-�_[�i��yUI������R�҆S��u�v9�Ԏ��� 1���Ʋ9fB� ��D\�����:����W?�QKƑ+�o9��Itr�$�i�_����"���L�5��3��嵨D�xO�0�����08<��f���{yDd�у�{,+������s�^���
���y�L�C�"����LD>7FV>�rV����?�A/n�ۘ����(0}
Tzy��(9��e*��̀���l�"Sq�l,߸�7���,��4I��Y�|y��.�V&M%�[,���e���"}��򨖊^�˷QA�A��)�'J�!c��tq�~��O��)Y�����"���<B��#�s��m�S�#~O�a��pv�E��r���-���}��J���;�t	v���p��¡#Iя�6�@�lvd�#�*1"ܖ�:��0��7K�T����)��hM�ː+�k�=��1�񵤏5�@[���N��;D'����p��9�v[�l���3a�)�.8!���DN�q30R�2��wf3\G�לH�;���W���B�޽�@S�3@%�B�gE�I�P�z����cXn6��'kԛp��0,��(H��OD���Xdͼ^n&�n&+�f��뱗�M���.��1��g'�U<��iwP�r�#M����a�g^��~���{)<a��`����b�>y.� �s���
�E�]��y�uA#�� ��vC��U�7;�$�����)���Z�������]�>5����BQ��@��S�e(%�yX�1v�49ME�5��L��	��$��`Wq��j=��u\�o�V�U�>�0�+R����B]s��a�-> �"k��"��z��6�F��J���B�ـ*K����WGK�Mw�-$���v=��9��58o��I&ѻ������K�M���`/Z��jf�#7o	����D6��4�H�떕� ��PYhb)ۮ�1��C��|�2_�sA���]��P��o� ��Bۯ�k�`�Љ��W�q������ #� �ܮ��3�
z��=�HLN��H�}���;I��0d��憊�=�J�N��� �=��A=<q�)�s�T����
|j�e)l笡G��b~���p�t�}$��v��y�$��	J�5�J hx��Jԁ8[6��ThP	�tP?�]t�HV�w��x�視���R��l�8�gv�5qQ��%!6z�Np����o1r`֞���GD�q�jZ(���L�r������B�.M��0i�c=��[�}���qjr���ʓ��t����jo�l/�m-P0���	n��Uk�!���*�.%G��M�l6k+Ш.�m�zm�>%��YL_$���E�ʠ�.�E4�b�h6Ѣ� w
��&Lү�{å����y�Por[ց��23t2+W����#j'�`:U�MJX����7.u�o��H��;,R�ǭ��-kE��lX:|��V	P�ݮ!cl�:�'�p}
���S;�S� b�⯥��L�Պ��9� m���3���c��_p��B���=��j�iȽ��mB8��FD*�;4Ez½�@�w3j�}s��3�֦Q݈Y.水a��7T|��as͡�˧ ��V�!�4<�"q(�7!-=�ٮ��St��z�TQ;٣�l��*X�L�}�&jl��\����n^�����x��L��FM.��N�����>\�X��Oܥ?}&�=����o-�¿�d���J��c�$�'Y8Y��!"R�{�k8��B>�W�^Ý���cg�R�X�ưVᙠy���*���;� b�����&�8�	��w=�o�Z(�� �����n?W�ƅ�H}a#A����C����@מӠ�QXgmv�c�̜?Ñ� a�r��6OϾա�ݛ�
���xKd��i��$٭�Q�K�TX�Ia����XU��<��e�	����,��2�!��pp��|k(������f��N��I���H���*4ǧ������X��٧A����rL����v���C9�O�:M��Ԋe�0�'�O? ����!��N�:�b��E�`8,ݥ��{w<�����c����C����d�o��]�+��Z��V����k��7<���5�����7~S�о3�H��sD��)N�G����|i�s�#�q%v#p#3u}ce��Z����v�� �dCL��b�i߹BYv�$�#*h{����fl�P���1V�I�(�j��8u���"�9�Ө}�p�_^d���'�]��
��s� N�3 ��K~���4P�D<��%G��(=�aI���ɷ�'Аw��h�\����c���:�V�/H��	��Q��xv�(6 4P�֟��LX"@�蚹���Q�p.d���=��L�z�5e�H�v��v�|���pf�k�Jx-���W2�rB�w�d!yI�l�/���[H� 3@� ��zPoG0[�Bkww����oI�fc {��y�i�Z��Q��C����g���Ϩ=$����'BS#�7=g�IY�`�Ѱ����1�S�Kk�Ǧ�<���/��iL�k_~j���4�o� �@�A�e���c�y�[#���H���w?=8�ڡ�E,�xN���|y�y:���u�)"��:i[ �S��Rr���i�t�O+X�ϙ)�R[q�!%�V�y �J�WͶ�"Wڍ�}��0�;�J3�W/�c*�h'2�u��$��m������������k!WK9P~=�Ȃj���aqP��/tE̅e�<,��bj����7fz���L��8%D��ߵ��d�W���%�!� APh��J$`! \���޷nϤ�]v�cP6��7�rtIc.	XƋZʹ�_�Ĝ�;�p�Iay��m�=��N5��eӥz��p2_iHӾ ]�ל�,�I@��"H�*J���F�uZϛI4mH?�� ��	Y~k�y��z��^��7�a��B�W��P�z�0=��f����M�Aۃ9�����?���F��s�"@߅�"wF&��DnÚ���g����w)~��۾�̋w&��O!�R�i�%^��&$:�$o����F��������w��ցU�K?��K}��u.��X",8����޴��/��8k.��8���Z�-ΟsZ���ܽ��tڨ�Np؉�L�u}��C�������휺�����q5��
3��Y�tҶwܩ"o\dS)ۆ�����d ��EV��LW���_����Dq�7Y�X��	`y*W���{�d d���\��˂.y;��j�IC@ϢL�y�V�F��P,�O���!�[�F����s<�H�s[�}I������]��'����Z��J��2ZM�G�RҖ4߬��Tm��o|	׽�V�I��G@ c> eD'bf���s,��5*.O;}ni&J�~�{[���=	�1����`�܆�	���}sl;Z��sE�r%�*�V�63��0��s����wV������JL��` ��1�?��ý�ֲ7�]P�9� �x a�h�%�q������(U�q���M���� MQ�OO������e�AnA)�GO�
J��7��[[h��ۻ���I<���+ �J�4L�~��a%�b��뤚-�hE�q�ڱ.K�i�I]�� ��m���9Ԋ���e��} �q��y���r^f=%��*�RUGO����Z�,/����CY�+��~M�T	3�Y�m�-�z������Ƒ�c��U�H��al�ɠ��֫��8G�R��Vz�tl�y����j��5��b��E,��i~�k[��Q1��x�c��oR{�B��n��[���v�Nqc��YlS�SL��*o~��c�n9��g^�#Z�D"o���@O��e�ܮba�Va�57�P��=��lӠ�4����
�Y���#�c���������h� ��>E��Tχ'��jc�Nf�U�iu<fT�5�W~^�@4 �V$&��^�j�(X�}-ѱ
'��]��n2��'��w��XI��3w�⓯��b<�E�)I}�"����������zE!�1�>d�Τ��|ڵ+9p ��o��l����1:�y��Rk��暄��<;�.�2�$>��!O���ECF�������8ŋ^����'a<�KP��niaaX3H�GU;�W�i�r&����_�aঊ�01�j�Η	z�-*2�J�x�h�A�q�Ƕqy��b���@��[)c?N��Ӑf3g@F�q�<�����Q2����۰y1M,�x�����6�ξ��b���$�v��s�:�}��E��JA1�t�*�ֻ�yQ"A�8��K�R��������KY3G:Հ��ںb�v.����D C$���q�¸���*eI��YT�!l����eLC6�P�|�rj4(\�'�b��vƜ�S(\�]OZ���Z��1��{�J��Z����X��d��w8�1,�1���D�4�,�)]�}h4�S|blTؗd�ϋ���Xtm�e�k��4o���"�a=!�z�/�s�׀��,��d�A����F� ��7d�Hͷ�����\�-k_nv�G�K්�l.>��~'�=������$�y���VG��hб�;u�j��	.Sɦ	&g97��M�B��~�S��[�d�_G�q��	�~�o�f�[8_�q{�����@�U��ҥ7�"����W
b��7%��c$�1���IR,��s��Q�D��<۝�h[�B�� P����0S�me�!�Cuf�D|q�J�,%{�F�9����#l��A����3��!@;V���ǳM_��"��+����ПP9��y���&���>�X�cL���	e� ��.ߎOS��:C���S�X�U뗖kl�I�!L)j�. Nǩ��R�	�����ۈ���+Vi���c�Q�g�B4���76#*X9Ꝃ}��) ��*)���.�⩰��3��).n������ c4�ɔ��4�LG���h�%G*/&4i���?Q��`�A`��L�-�BfC��bR�鼂k%ҙ��cҮ��n����]|<������2\�� V�I�~�"p��)�c�m�"ODL{�T	�ʎ�F�s������fA�6N���+U�~�m��q��)]��0����ɗ[�c�:�_���۸��Q�c¦]�k�yi��_{Ζ�E�S��D4Z���/�f.��Ҿ��f#���㟩l�ݽ4�+�02B�DM��R5{�ZV&p}�\��po��EѾ<�$?
̂���?������aGw��?Ql��:�W�!#�(��y�y�_�� ����k��SV�Xz�.�� U�I3FN?��էU�@=���9ɪt
N�+<0|�k�gFkj�a�������|�O�eJ��^VN4@q����v�[5)�C���m`E� ;ҽǺ%���Bn�Lk��������f������ ���f+X�����,P�uk,G	�_0����<��_��/�Xe垵ILN��.�;d9A6Z��I��'��9��T 1���䴴�/��Vv����{�m�)�#� �n�%.�}O���cN�{���&�t&�1���z-���Y}r�����C6\��u�!o[A�E!V*��o��t�
B?��B{��0Ɗ[�\DC=�HZi�_(�+�{������z&����p�"56�z郠���� ꁎ��M�G�MDd��\1��J���걻�Ⱥ�rz�,��I�2hަ`
��ӝϢϥ�Al��J=H.Q�|XZkH�H���I����������0Hx��̃�oLe��5rZuM�nE�w0�@�q���2 CvaЙ����<��<!rۉYux�Q}�P@��qzO����������莁�|��߿���; �Z�<h���� 1U3�Q�� ��al�n
E�j�jt��>������$��{I�މ1�kh�\���+���0GL�N��~Ls.R_��9��9���`O�9�)}D���d���X�6�c�%�o���D�޺��w48����f�Az���sI&�p�/�(�רa��7%�@}��=V@PrYQpY�g��@�Zag��y�����؇w���X)��yD�tE��jjj��h|��|jo�1��PM�~�S�s����H��78��oF�m��(����$zo��n���t4�k�����팚�h��!/5���c�<4�cG6ZFR��?�5���y��c�^�=H��vFK���r�=��>�4��:|�C/��,\��T~�E�Ω��oi�#��E��j��N�[#2�C��Y�)��"a6����X���M^#pM��i���O��'�2"ԭ���B��毌���vS��J^+:�t�P~7"�B�����xM�.�&TB*%CPUJ��,�t5o*���,�nS�����G�At���Q����8�*�s�Oi �9C��<�̉�|{��Ԁ�P��T>�%���f���335���x�w��
�:
Z䡴O�N�i�vT^�ܕXkAX�ȵ�����%0�:�4��	�l�-k���D�������C�L͞huk��B�[��0���E��K��������E(��/&
�-&"��P��
�����;~�q�	H���2՞o����mk��ixQ��	��јA4b^;7O�nJ��~ƺ��8�$,��~�x��$�i%���qC��1 <O��C;��(�ڑ�e�^=�]f��>�ohz齀�;j��6~�l��DF�}��M�t�·*�؛������,%=�e$]b�?M�� K\���[�!��o��p��%���HD��8}D>��K@ɿ��MEHv�$2�.�T%�옣6����L6�(k���;��=�ئ�x��v}���ͅW5�G��c0hg�T�&�|dF�������"(�|�p�ts�$���?�J���W�}��)X˥�6�y�1e=~?/)7ȗ�&vI�2�`	ˆ|z"�8O����->��R8e�n�w�+SvWt�|[�"s,��n�����s-mCY�Q�҈���a��7d7f�#G���	�I��%���{���P|G�.�z�q�����/@^�n�\�~l<c�$q�o��D�Ea[ןҿ���� W�����w|�h��4uS������ u�����c(�\j��O�w"<�K͝Q�*���D��L$�&�0�Ņe���D�)q9��)�=e 0�2��>	B�.�:�Ud�7,���+'Z �d���� ��	�<	cu�0U|\79J�}�c�h��"E��n�X(WN~WK1�������@:�����Y|����H���B�b�X��6m���dN(.0R���S�"G�����fq�	4>����� $����p*<3��G�G�Tm���=z�r���K��@/xf��.������Ȍ{N:m�F씜����� 8_��w�"��c����p��	����4q�o����/�=��[Wv�͞&}�!J���M�f�SN��@�w0��mh������a��M��b��q�j���t5�4L��'2�O
�ł���LKd�D/�i@� ���孋�:c��u�:�����*粍�mz�{'0a%Q���m������u���ujf����s� Y�)M-k
�������O��ICۧk���j*������):GNV��EA9�_��7�$��2��Ec�1.�ϯ~�DC�*��t�o'���X
K붳;����>`���9��$��C����Ҽ�ޖ���@�;�I�s�>K%�Ϙ��*�ٷ��K�<��q��ݲ-���3�p{C+p��i߻�!|��=$' 7=N�rM�o��{Ƥ�c�2>e����������`�Tح1�֍�s����!4�̠�bF���7KP��\����Vbߘ����+1sλ��*1���&���D��!��iK�B0��`�Eb����K���x��{wg���hͬϞ¾��P�x�b�����Y�6^�¿&��d]���ę��	B�	`�T��ؚ��Z�Hֳd\H!������ֺ����hJ'*�):g;��9��	2+Lf!v�p�������7�Z��\�hA��<'8%̣7�'�5i)[��