��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ��(w����E��}�U.��K0��m�A�x�����m]�ǟ�������"m81T�A�q��z���7��M����~�`�]����9�Q��qۘ�C��
�'�//T!�ѾbA���sq�]��[����A9���:��+�<��s�A<����?����C��A�5��i�NV�V}�������X�R�R�=���\H�2ŝ�`tw��	��v4(BT�����:F�Sݼ%�+�=�1a�M���ދZ��q�7�/K���:	��&�_�V�V!.6?(S��o=��m�4��X3ϥ	�6��ĸ�����&����2h�� �la`��<3ۈ�lb+	���=�N�z�RDn���t�Q��R� %�HN-*o�}/�p*#��Ƒ��|9���8�4OD����x���	3�j�ƬR*yJ����U��>����t�F�rq�P�V ���y�r�v%}���bK���>����?�<���׆�-7�:�/2��l� �x�UE�৵�R �#u���f�(Lup4��7(��6���v�:��U-�3	��,
W�sU�)���F�!ֶ��Ql���Q6��Bv�19��ͥ�f9��O���L��2Y�u v��D���0�}��d����f�2�KËa7��H�mN�`��z���u�C�N�`?��o	�96��`��� ��EX	���T��.�Cu��m0� �>��[����A�xp�5��֗�����'���U�;��ݒܠ�_����pEeOf�3f��(���B	4
�R"|��X���^����ɉ�f}A�g�!��W%�4� :]�^�%'2�����߼Kzi�`n�*��"b�l-4�d�����#��ȍ
a�+����ywR��P�r�c�?�y��4�ײ��|>H���2axz�ڦ������%�v���8�t�%�zXJ�c��}6�&�WǱ�:�矅#p�����|�׌:D��"��#~�8����KE���FF1W���^R�R���1�����@{�	ct�N�C"��p��n���B�Y3|`Vd��������ψdE1�Hץ97.9GW�.����� E�y�V��'�Lz�UE!�	�7Up���9��&�ck��bQ��r]ʲ~d��y������_4N�;wd� �bz!?�@j~�v���)*��xh�*��^��N{��{�f�aa�^A����dh�{�q�����^̮�^���q�����k�Ǡl��[� io;:y�����5�W�҉l���/i�]�E��{^\o�!2Då��
������M�1ũ;C��q7Dc��d(�'�������f�r��37�#\2��c"먎�*��=X��̓A�����E��ݢQ}NV�@��W��8��Um^�R�>��?�[�'�����	�#�H��ҁ։�����+�LB�3���v-Jf��|p8����|���[A����OU�[IU,6�ȼ3f��\�7���`÷�(:=}������y�6�?]�3��a=}a@����ZF��J�\�ApD8��8�{�_9��~Ʈ�M$z����Ǡ�R�G�( *��sg�~f�A`74�(�D;~8��p�o�����S�921�l�\��8��-��7�����]\�8��y���+ݯq��7��	U�"Q���w�m	J�ii����#��H�$�F@�"� hj� �ߔ��]�/���uJ N`S�c \��[�g/#���KI�38B%چ�	�.�;�Rc���WHC�O,~�vz�<��.�hebT�1�q�"�F�mI��㶙RX��[U �o���o~��H�y���浳o�~e*Q�����q�<��t��s�����H*&��TBӑ��0F�|+"!��2�n�P`������);n�lU��x�s0�<
��G�Vu��C���UD��6�Wcb�
D�!����{��?tr%�d���6e܂���گ�X.9��&	��XH��n��i3�>����(�:�2�\�%���W2_rL�������^��-�D�ϯ^�Oa���ɚ�푙���$�k�$��.��i��0p���e_���)�;8u�E���3d��E]��я�'�11�
"b/zލ�6a���O�#����ug���;p�h#F��V�)��N�=0��v�Q��aQ���)=ݻ}����ګ����j��߂E2k���e��˨Y��C�_@�-�����0C����)�.�.��h�_�"qK�h%�n�ab��3'r�O �D��{]�/:�u�0�l�ȑ���^>)G?���lV��HZ�V�U6���LՌ� r�1E�s0���`��jJ���tRⅵ���{PD�A�]�R��{�Gx�^�����yk�wm�?��@��K'�	j��Ź���񝽫�/R�j
��CM%�}j�1Vg� � J�a"''�#&C�]++֞T{TW��1���x�j�
7��w�J���I� M���o����Zj����ʡ�0t0�i?&0�䙆0Q�����
�Xn�W�LH6T_��@�3����.T.A��8���{!9d����4Pu���p�}(��9Ȇa�t6�P}�
�H֋P���&�E�t�PB��J�i����&pL�E5�}��*��EB`۩�G����gO��́q0[� ��IEd1�b7�Ia��=6�.��Q�$�Zx�jڂ�v�Ѫu��;�����SqK5��'\7��D�r:�̪hf���FBT��9�(,�dr�ٽR�%�������:,4�'0�Z�$�kC�)��)[z+�������T�U�&�=ρ�?��F��� �e�5Ag�ndIv��[�Y��?��\*m����QĴ�*���Q�As؛���O���o�`�=�{E��S��B��Roh���SpC��R���b�$���	ϓ
P���^h�^����CM���ʜǠ��"FV�G��b�A��Z]�?a�l�rE;^z�LV4;��K�?��Mx�0��DV����Ϋ����W����l���1�I,����_��:�>Y�>��)����;�V}8a�+��S�7�J�?'u�,��"9��i�*.y�ښ�gpx��'�)X+�T�kҁ$k�i�2��
�ѧ}u����f���C4Z}i&���F�|�<���*�[1�lֲ���&Kr�Hi&-d�p�5M9R��v�U����+��ɞ^9F���������m�<���;��=���7�{[�@Y��pOh��63r��V�D�uK�	FmK����l5"�J����`��?���M2*!r�V�V�G�Z��
��n�;�$@c� ��j1�E0˕���,��x�U:{h^�dY�L%�@"E�@�Pa�'l�:�AJ���4V�c��4 �O��Jz�;i�:<��cV���!�&J.�a���r��p�&��	����C�8w6����L�{��R9@LN:<�`�Xl��8�k���p4�-���1��e�2`Қz��r��)v�,	��̢��TEX�.֍�a3wҒN�-�y<��urH��x�Z�k�(�gQ4��6ڜ#?��:����6_b��v��l�`��z�A����YWfm�ՄbF�
����皀�yD����w6�q �acEՑ��X�~�$2��1�Џ,�7���j,j������O�ϳW��}u�@F��� ��7u�|�q�*S%����R��U��dܶ��a�(�|��*�+'�r�G�V�8+�i[����.%����r2XA�L�N�[]9&�R(��L&-�4{�^��Q����4��\>8��OW������ڈJi���$�jФ)�����Q��i���w/s�r�P:�+l�	��OFU�߻�+1P	�:�`���gQP���Yλ��RV�%+m ϴf���:H;�/i��BFL���"�_cf���NE�Y]qO������������%�mK��D��!�e��+@�;��
�yRTuu7��sr@^^�C�}�fAp;s���)�D���<�	rE�W�`g*L���?#)�w~K�Y�N¾^��eRȔt�����׮��\"Kk��à�ќA��K��qd���I�?�@�=gz̊s��DKB5��c�����B��p>C�'��Ff�rs�ɤ�_P������ L%�XÔ�"\�|�F�h˦f��,�ڢ[��<��r�5���/~�C{V�0��6޲To�a)�I��x4�&㮹���M��Eձ\g���L��`��������H*?���ޫ�}�E!�����Oe4b�-��z�R�T��~c�>���l[ϻ��&�F��f'h�}&[Z��+�r1�
��:�k]�՟t�z��@�x̆���p��:�Q�)i�n�x�ڝ�7���[��W`.w�ɺ6�&�6H�����SM٨ÁL6@\M�Zt�A]ZyP�,�F��}+wcE����Ym����t���G�aGpև��=�nl\��A �M��J�x��'n������;�N�+6�l��d{���D��uu�@@��m���a�R�p�����O�`
�T0��������J��f��7��%��=���xQp����b�C�,A��wG�h��Pin�r;����0��M�8E,A��z�Ҷ�Le�a�;Ҏ������7q.�����SPb��K�
?��LQ�7��U�^@O9��� �"D���kW_�hy�����L����;��/��~��f�YS������x���m�^�(P�[���h�����Ƣ�սc掠��E!�6F�*a�p�44+��`�w����Fj%-BD0�ZB��A)��	�#�~�~��GòUK�].!1��{����=�{��AO	%tzl�1D���K8�_��Xx3ڪ[�9c��Pm���#�]�I�K�i��\�-K(�����"V�"���&&�v��kLR%�П�������F�zLu�+�Pu��]�����WJ;�5�C{��{�_pb��!�,Y~]�l��v��O�����4{����Ӂ�n�3�tO��1�f��#�{�܈9�0sk5���S>t�h�vQKW��$_^���4���}2�G"I�����w���<�����Խ$̱�ü�����	K�J���iq��䩍��ߞ]k�v�Na�|�%wJ^h����|�{�Y�F�s���ʂ�L�)U��\덤��c�Q��+���� ��L�h��E�,�K���F;Q�/X�O�s���JB���<�_�;y��T<>Nn=��/�w2߈Z���Mj�Hrt.9p��S,��Ӣ� ������%���v��Z�)���,��H׿��}�CՖE�=+ �am�P ��i��<��a��k|^�e�G�{�k
�c�2��6?O`���FfH�ա0�dF$���4��J�De!y�W#G��\�rZ�ʁc����_ �WZs�0���h4t�-�1�i]b�x�fg��Zody������ �$$�=+��3:3��ӲNeF�쥑��HWc�zs����k폳�5���#�a#K��E\o����V"iWL�B� ȇ'c���j�>�+�v��^�Ć�-�Q�H¯���Ul���/�2�/+����諈ӳJA�Зρ��*��:�Anr���`V���~k��,�ń�;���x��[2��t��kg���{����oÒ
u�RCGLKu6X��VX�LԐ�H�����>Tt3���f��1�?zq�l����{Kc��d�-Ԇ��W��Ӻe�i�u��2Y8�lQ���]�oV�Kk�v�#2�_U �C�'���EzXM--�=,��(u�́�{J����`����|� ��R'�Ь�ax�^����o��#��R��(�1j���c2�)�
5�9H^�����_s�e9�z�z�Vݏ�
B�h�Y>^\#�����UKn�|�K������ t�2��+�O���ߵ	�4d6�նn{��Z��}��J��-
*_f�ۋ����Į��H�a�>
��[�,�A�[�t��ih^��Qן����)bo�.3#F�w�4�o�z���(V��Wîc�V���.�����U�;JU8b�B�T��c� ��M���w���z��8
�]�u0��������͆�o4z�;�P���2a����7J��?�~�S#J���.F����6{+��Zg(��Ŷ`�94�k�/�Z6��	t|:���_X���NC-�� �^@���,��}�ܮ���T\,��!��s��:P��-Zp���؃���i	p׾�!�X^{^���"������K(�WYut���ax�ϵz������v&�#`b�'���
ٟ$�>��6E��<	�k����y�B�'��ԉm�W>C�|�?��^ߜ�j���qZ�-H����o�U�-�i��Bā��`a����B��0�Xֲ�	v>�޷�߈�k:sB5(0
0������z��u����8�<�Cf��eG�^���JcVM�:]��V��_�;Ø���..�7�ލ��n#��а��CMZf#�q���Q�T?Б$)dމ\���B9��Oa�B�P�Q7��N�V:��K�r���R���`n���щI��k ,� �,؉�W3���!͆nV0Ė���I/�|�c�h��<E4ޜ$�����A��F������@���*��:����w�T]@�n�9S_+���_�w>�������/�[�o)�!�q<���$��(3��~��G�f�w������_�\5�H��w��.#�g�N1�0Y&ځ��UYCr~A���.��d���-իצ>yƖ ހ%���V3��H��\�?�`�D1Ӿ�P��9�y ��:���D��v�`rFdo���d���,���ȋ�W9<�X�ߢ�� �]���#��P��WߒZ��5 e���T���J�M0��]�ٮ���jpz=���
p��k!�\��!��N
g(�tB���uç�+�b]�C\~H5ډN�N=����r���$�r���5�`i���#/86��<��UHDY�U�`P������O��4tr�|�X�%3�����mWGĞ�ě�>��؁0޵��o�3��)�պ�̂����(��M��+�]95`����ͭ�������~gBP<$� uf9y����WQ�= u8�o6�T'ܴ;��HU��������z<�?vl� �Z���bS��d ��~�	Hj���a������ j��BC�!)nGm�#��g&NJO4�u�����vu�X-�F{������O�O�8���ےw��御���)�a��f�m�4��3�'3�mī·Yu�E������7��[��֋~�v=���N��4�a���S��hR���@{��<{f�K��1\"��p.:X� 	�q�|/�����i8��@����H�1�� הX�bӒsp��u�>9�N�{[�m ,ͧ1��Okh�8�{�Ç���VLl�&J��qO�+���\v���j�n'��\h&���$�Ǵ���o�R]HA K>�3�`tⷙ*��?ˬbD�9z8},R������G�8Jp\�������Rre��d����=ҔW���L���p^� �4%"g5��a�_����T�H�3R���֯�:�	��G0t?�X�SH���Z�4���w���2�8�o4��������}q��M��L�/�-k�`*�	�Pt!�$h��-\��ѯ���&.�1V�)Ż��m��/��NTy�A�E�!^��ϻ���/���!~��-��`�V���=I����w�w��#x�?�N��0�w%Vڴfz�F\��[�,�
ۖ������q�펿���ν��P9��l�����E�r�zj�a��X©�_��Ja�I�(�,��C��T�!�����/`D�eN4ܝl�%)^T�YB���[kQ��ǅg���Y�/5X��0�@QD�tʁ-��Ƭk���+�}�rg$��4(g��u"������91�g�I��PZ����.$�����k�_o:���'X��2���+7�~�' �������w�$H�c�8�Q��gH9)���M�!���ֲźW�l!��{M��Un��M�G���uUi�z_ `�fB��C�`��wP��],�p=������ɧ�O��eDI/�19�z�B���߳jõVDE�۹�:�crH>,E�H��0��`,?��{���=Ox��'\�����Z\LA�{��(�S?��C�]*�ԫ�!_�n�A�_y��gt���ˣ?�ש�8�($����a�&;�"�+�a��*�n�X�w�(j*U,0<����'�k� �q�{p}��|�����!m G׬׃K�ˉ�ؼ��t��k*��9+ѿ=i�s5^������|���|����b���5�����{jY���ğ�-�#E�S䭴���Ǳ�4M�0)��2�:��@�����w�E���b��H6AW��1uL���x�F��@�= �G|.���ī@Z�Z�x0�<���?��B/[Zɤ���曌_�Φ�����fM6�K��/�qH���\��2bx"f#���X�(V� 5���Uȭ;á�u����SF`u�9+V��� ��|%f(�
4q=�U��༴���u��Rk"yi�`E��`��^�J�<�q�s��#�D�5�ӽ6�2bC� ��L�rըV�$K�{�O)��a^�� ��PR3�sݳ��Ǝc͝�+4j��\%JԶ<���=5^��p��2Ll�{r�0��f�I:m ܫ��
^�d�	J�A`c.�}����:C��?��_�$ϙ�0�l�X�L��kwZH��ߋ�7� f5Rt&�!-a�0�xOj�yW�J']�L2��.� �pӨv-5=�wM�l�£���کM>=C#(8�Ө
�1���l�b��
kpŝ���'��gi���h�� X�b�H7�l��Y��������j�̡��:)Yyx�5t6���9���S~���
���'�H!���e\���=����!D�����,���4�U�>a&���q/N?4��X��C�4=�� Et�m�E���͕���j�����%�A�g���E+*�e�e[�&!S���OQ��a_p9b	V�1L�Pዽ֔y��s�Ui�5.Ç��K5����Uۺ�m���� ��Ci���V�kCv��A���u�1�E�(�� �g�x69/�ԋ�vT�F�!�%�� ���iR�cF��Q�����M������]Z���vi�KA�H+�����*�p���+~��=D$O�:{�x�ܿ�R�M���z�3��%�����X��
��U2�v�oo��(����=����D��pNoFp��zM��}S�48�}����ч��<�y^�H��|� j��to�&X���:1��"�*O����@LM7�Bvf�*��A�D���|2(��o�S!ҹ�0������Y��w����L�9���v��o���u�e��]Cˠ��5�9���}D���E�QS����7Qg띤ͭ����;����em1 4�S��������l��bSݼ�l6؁Â���ۓS��w%�����P��uo`��Gn���7�0�^x*n}P!�8'�:�cm�ՆR.pJ�n��c�4��:r�rb�]�au��_L9���2#B[�ʀ����`�Cj{�~jZqD�W��º�����;D+m��,	����I+��S�js�k���ɝ��dB�i'�V^����O�;�"Q騯۟a}$^l+��<��������X�8C�_�V���P��t �LY�6#q���k��o(�V���?�i��x&���k�]�`rR,���{T��a`Y����oL����h����76�=g�����4�˽F"ONke�6y��Z�����=�XLtF�t�v���^�(�%�wW�����-֌^����2$�"W��$JR��h�.��x���_1��y�J"����u&�r5�c���E�Cc�����`f��s]4�V.��˯Q�@�f�6
F�l���+�튩ݵ��t�[�08cZ��\ɪRfc����R���^RFJz��NP�����������V+"�B>[_/6��j֬ ����?"�u�p�<e���/R�ί�n&T;�:����G���.�j]�������E�ɷx�v�b�?5�ˋ����\L�-ݥ��b���9�S3I�+#�=U(�D]�d��4��qmnYj��TXʜ#V��w�u1��z5��x'�j<�*����e�{����Ӿ�Y.�>�)&:�!~T/ޕ��-�˦��(�6xS��Iz� 4P����I[>�w�l��N6
&Xs8X��9h�Ta�s������7.�ͦ�}�c;��%FF^���1�yE���l�
6����K	���T:ܟ3��Ə����-/�����o��D���,��u�4V��CC�=��4,16���o��ڭ�mr��"�#�*2~m�|��n�ԝ���Y�q���ԕ�s��Z�������h�Q�v|fh���GH8{�B}#q��
�����^���%0���Wl�tZS��V���H<~�jq������[�k����,K�wKw��B}��J1ϱ�:�0�y��{df�V�}��ʞ$�)��0�v��V� y`E�>���DS仯(������w@�� �jʮ�u9��~i'�Ͳ�I�J95�^
�F�=g�l�x�ո+�(:�Mj���1�u����^��?6�H�e�~B�~R)�7Y�za�ĭZ$& /Q���fB���B�c�t8+_n8T��zK�)'�7�PJ��ę�G�*h����_�lND�`���6�+�'���Bs5X$�9�2aG���[J�0RZ��C�nB���]^�t���DN��x�f8JBT:��߈=����������@�W'M��F��ٚ��Z�����cAU�G�L��4�I����**��!�M��M9���u�D�Tm��oK=��3��+�U��?�C�Q"�'ڍ�ql���/r[>i1�=�0u�[;��c�jE"�#���+W�V%��O���3"�ٷr����p�~�@����\��H�S��²m��xmk��ѦԜ ����=a��I�J�s���vR.�S擂�^��x�����ҭKyȾ-b��������������w��t�?�|�O1֤b�+����/Y�����];8N#�L�H���領�şd �	��ե���p��v�OU�;�K���U��ƎٌQg�9���H�����Cٞ=�}N���@;ڀ���ȻJ��1�pY�,b��O���4�X�C��?����
P�?��Ϭ��]��`��B�I@�[RO����&c���9��Y�0������v�QC>3+��YR��]&QMY{����D�0��~�`4��3;}�o�!��Ut�(���n� 5�����W��k=�I�0�vr�ڥʠ���+(���Q�%��sZ�uL6&Y�:
��G�Vv�০6�}
�� �D���˸��,�����x��O��%O���,6�5����7O͵��@lp(�>�ݲӷ~5>�1փhI��e����O���'ٺ��ZY�	�H�ā�J�D�p�Ics�n�M�2���Ex�;\0�􉴩���"I�?�"�� ��
v���#����?g�1� k�=�:-��l�������<X���M����`��!��� �y4U���hU�ej�/+���0�z�Ǖ�˒�O��o�'Ef��Ax	Q�����Ym�*��Y��09����R��}��e��}nz���F�ȷ�e&������N��>�e�#��,��L|Y&r!W:U*t�����.Q����C@h­��&Kq�.ۀ�]�R�#Ȼ;����ça�$�h8�����)������0:F����e���yC�@9&Ë�X�ju�y���.����n�8y$R�"tpU�ô��ۉ1��z����'1ᨍ]�sK�l��aq^�as��v1���7�nVD�e��Y�S�gdr�D1kz;/�11r�/���_�3�l�$�]�����]����t�'��7Uш�wˇ��J���R%�VS;Z�e/{e�N�9}+����=C���%j2�0m"A"��fԡ�c�;5f�G�x����Ui9�X�	n��^��d��Kn��^��avm̋g���EF����)�<�g�l��vVUze�}i炂H<ByW����s��U��>Q�ܪ�ebη+���.��H�w��օ�u�pJ%G(*�ɦ����/��.a_��'�2��������5ώ�s�zvG��M��2������~ٕ�@����=B�|/Y�BK4sk_��˥��'tO^P�%O���TX$}���~#vJS,جuOц��\��-�'�k#�֞;a7��I�r��!��C�����,�����[�
9�$pc���� �������N�ڗy��ʹ��|�d�H~�☻*z䦚�㟘w�^_12E�+:����Q6�LL��-r�7i�� �_�D�����ꇸ���H����Q�Ld<��-#S��O����y�;�\iXKQ�K�+�~Bs['D��#�%gCZ|�bC�1�K�]������M�;4�v�
HL�+o4
dG����'CN@N3yN6�#��5(��<MmEv�����:�p;�P<��edi�-�c)��t8E���xMO��P������򿿋���p�*ЏS=M;�Y��M�Jʉj��&�qi�%�Bg�3:���z�Q�cǙY�G"md������d"dDg�-"#7`mC���E/���Q��I>2y!��c��չ�u���ۤ�$�]GI���T	O���w.�z�.�����Ҟ(u��[)�>�$�\��	��W3�l�z��qz�,�T������ QzY��v�v"y"Vb� ��жS�z`x���i��T�L7bf���7wJc�B�Ayd����c�n8���������ϕ|�]��2�X.��wr���_��=~�c�Ɲm��@=��[�`� 0����xH-�c	�����-��F�+{ؤ�C7X��sP�8� T3(�ia��xt>�rN��ҢG �Zm e"r���U�ĄcU�9�J����_sn����W7�����j��WlG���fj�i!��u��Il�\�V�M�m��	m�'XNr.M/Dvƨ�]�xa�I����j�*Έ�U��4��g��`�W�f^�c��'߹?�`g��R�ܼ!w%�k˯��M��=�,1��3�T��7������M��s�4a��R��Š9��BA�^ު�xX���!Gj�������pI�Oj��#��[e�^=��TG��G�$\�*
�|uB���v�R*�3���xWO��+U�0��Aʽ��M�;=)�)ү�ZLB Aj�7�����bV�1����$�\�ج�^���v5P"D�`5*��C]�2��Qi$4��n�^򁧻�P�������!�|k��̲���\$"ᩀ1����&�U���/�*hG�{�yE���pŷ!�$�_H��N��:s���z	|>���e��18��dW��!6_���S������K2�ҧ���z�-�#�;�XT|UQ�V@4Mۉmu����K���W|��;yT�P/E.^*~/�S#
GޠN��P9A���l�jb&���Q�UfɅJU8����3�Ej?�.Xih"�<I�4m@���R���\�*��AK�0��*��u��� nG�&?%����.Z�9��`(��z�]M�;6qM�lb�dD�����8V����'�������n�A�r�=L���J��t��*)3g�2��P~{�����Ĕ����Cla�m�1"Wƌg|˭-L����S&���+��w;ȍC<f)����g0��u��լ�*tg� ���$}�ݧ5�`����F��W(���,q�?�;�x�4���c�M�.7�|^�hB�g�i(*yQ��D�i���#�8� �0`W��3k�jF�3���ij�as�����{;\.z����A�$��W٪�ci����oJh�f/$8^]yػ����M�]��hɇùw�����x����;EiW���T���𔴜��Y14 �RfU\q��IdҘ���0�R�2:�@�I���<50������ ���t��Nw�84n�����v�~���n�&�����iڒ�����e�J�k�z�J�]�̆�C`MU|O�"����q�/.؂
`�\�ܤex����>J�xE�V��ݼ��,�gY�-�/�:t�(�p����x�S���e'޸�"F%�^��Bc1k&A����焇r�9��g�-�L 7(�X�����V�R��R��TL�8��5�&�L���;�n�v�4�1����6�Fѡ����0��b\B����3K��F�,��X03ޘ����QYz�-�N��sCp[���s�\��˲uxAu�G"5�K&�i�d��
���喒���LQ-_C��59ފ̇o�n{�X��i��j�Z�p�\RIә�Gl��1�c[�;���,��}����͑�'M��.��B�ud��~��=�4
���DM�ׁpGb9vjk��[�wM'*p�i��W_S�U�z�ȿ"V|�����EE�B�Lɶ�gi6����k��6[qB{2��}~,QR��S�m���[�9����TR��9I��U��:�Z���a�8+i6BЄ��WE��DAV�U�� `�B��Mk��֡c$}����GΩ���zVa�^&9�]��Q��ʕ�Qb���N��e+�/�v1̆��
�@�������l��)��nR@�o���ݘ	����ahՏH$��kHnI"���g��%���:X�*)Mx��*�6-ї3m�DOn_%GD�N�ݏ��u�!�66�č��-�J��L�r&��9��U�zC����M�;$s���dqcR�{�M\���#��͛��n;2wL}�t���7ܯ��|@69���u�/ˠX~[Tf_�} Ȟ�-�Bt�D�����GɁ��n��v-5�יy�+�);4ei�iM9m;�H��q��7��ӄ��1�L��4�i~�:#+���A��=,����"Iy��[��������.��7W�6��~t:����P�q��h��q�+Ħ��g@��Eǋ��{�nK�Y�ͬ����8�T��������^z�>��=��8p��Ww�
9�m�?w��_x	��=���uo�
Z`�hi����l����2<����$�}(��ߛ���z�E�$rX ����}�=��31צ��\&X�(%r�IU��(�2S��B�V�m��W���un���O�a)c��S1e� �ֱ����;bhi��Z����ħ%�Ο�=&���@�M�S�Y��qמn	ğ=$L�m���L]����Kaz�n�y|x�--���؊����9���#F��\�������ܬ|�Hc ��K�/K��1Q�������I���d���:(���;�.���M:#T=�(]�"D���$M2PEg[�.<a{��l=��5�$(E��F�g=��r>��ZL��f/�$�𭰭���Q[l�|�O���!,Q��V���9��D��x���,�.��~W���&e��[��(WD��;��:A�bpQ�3�a�I�c�:�[:���{u���$���3N��<zYN���&����r��%G"ihnjA�{���N� ,x:�҅����;:���Ig,(�%Qf�c�=tFJQ`QG_�M��6cS�?���J�}� cTLm�bpTg�s��J�T��̺���ϨRN���ӱ�9�Б���]�R%C�����_�	�&��H�,�n��񏉒�|��,Ӗ���)F�D#�M�B�Mix���J�����D�-����"�w�L9��Ҏ>]5ԑQy�]؈�3R���g��̶�˳�N���9�=5(ܱ��$M�\ɳ��_��6�Y�Il���vF�r8x�:����_k������G�Z���f�!�bx���X��Ϝ��SCӴ�����",���٩�d�~���H��30��INE��Bst4�����)��<.Ɓ8�,����z�,�■n(�tAvfXn��j�CAg���M���@餯k�Z:L�^g��W��b��$�Q�䄡�8����F��v���%k��T|F����3y��Gn��t8lf�.K�Umw;�_��,�1j���9 Z*�|!�#t�n`�$.o�`��׼�����W�jhs�������>�"{L^�oC&Q���-�O�u��5�x���80�j^�8~Q��Q!�?��@$��c��)�F�D^e��}K=��]�ROC�S�/HHWd!��订H�7S-/ɓ,�[��kFO��	ZmAA��F���UB�5�Ղ�􋀈�A�E�]����|ȟJb�~?����"��K}4��9�Ӳ��f���z��$�<��e�uk���JIv������!�C@5P��n�Nf��=2������]�HVn*�	�=Y�Є�-NZ �ε�Wo3hj�3q�B��=^m������5��%k�u�D����1��L��*R�'�_֢�b��c,a��m��x�K�!�a��K���v:^0,Wѱ*��]�w!I���xO�!x��U�,����Ґ�A�W��t�m�9Ԗ5zm���N��\�%�x0�ȓ\6�0�<f$5f,	6ld���*����D���0����(�7��Y�]����SB��v�k�Jn�3Z��X%�j�C�޸Ք�UԴ��M�AŚ�,��֑�;d��)uj�"A-y�RyA:\��	靊�V�g����A܄$�轲��������W�H�#Nr���f�Ia�Ny���@2H(��b�� R�M�N��+nc���`T�E)b�ߡ���Ś�*���
v�s��)�I�����l �Uށ#���V����čW܀}�qp��Csf�&�b����%���<�2�(@o�YCDu�ձ�����*��"�~�H�� �_�,;#Wu;�֪N{%�	&>cmQ��!]N}'��e�j���|�]I8T�<�E����4�賖��|^%�	�������%T�7$T��F�]���g���JF6;-��@5#וS'z���H�%�F��k��3�Y��'�N�Ov�������r����Y��7n~�ĭ��T6	�����>i}Pc����Q��ߒ���&���#*��	���)�ڊ6�P�k��M����G�t�	6�^�bC��"ܛ�(	#M���nLF�����`��
HQ�R���X۾�����nxi��R�`m�fz�v)�T��*�UZ��b��V:�}�#�[9F�Bę��:IH���_�����0����WZP�)�� ��J��bY��'�f�J��o���NA��$>BZ80�?�`.���0�B\%�z��%jDC�;��`�&���4�*�h�	�W?p���sA;�(M����Z�:���0�,����M��ܕH�+�y8�S���3�6+C�|I��ȷn�7��C����~�-�p�����H��8a�5|R����JE �X��yז�i��[O��X���[1mZ�b���zEٰI�U��4|�L�Kj1�g��� b{Us���?���
��_�5����kgo�D��u�vV�����`)
�¥E�{����7nu�Jj�B�K�0��I������gZ;5^,�:wn��7B�J�h��j�����Ц�m:�dF;j��\QU�"��iyh}���a�צm`}p��Zl�u�غ��|�?@���H��(_'G^�	p?=V��%�v�H �$�����_;���g�(Ҙ�T�Z{�滛��m?�����Oϭ.�wl��Q^�s�l�G���y��1�����*�g��,}rՋ-����Q�x�����{��(.L:�.����{9}z��&��g�~1�Vp8�!�>ݺ��Cj�۾�'EMZc���� ���X�a���F7r^#�;�n�����Uqy4�/��7hqL8����EF� ��C��񘩪�T�]*�Q~�L�fB~ F�M�xߣ��m{ur��ؠo)�絘���;�m$ݶzo�0)���5L+'0��XIە��cnq��o��A�>	T�%~m9�B27�Q�,Q�T�Y�7�懌����S�#��L֖tZ�x���������v���_D;��̀�OUVHՃ�P�L.s�_��p���w�����Y3w�D�jƭܤٿR
��
Ä:�յ��C.{s".�+�𣊕�Y�C��4��p�����%���$�HCr�Tm*ǢO��@$�X��q�9�mF�v��СC���q&v�N�w�@�2ȉv��i����C����i���\/�,�x����<��HR�q�*���$]g*1%�bAխ����n^�Z�ܩ-�j��L<�(aED.�yQ��d���Q>�#X���n�y ��Sr-]��H�"8Ù
4��H{�is���VWe^BMCF|��gb���?�_����܂k��?HNU�[���ck��X7gɗx���P�X֬]01�q[`�B;{Y���ř�[+OFgj�C#��\'���0�)drI]�[���ұ�#�kG(Ojt�����X��5�2�Bb��T�� �
.��}I���S�Ȉ�0vǷ�>�T
���t_���ge�����g���/,3&r��f��yt�<J=�k����~���u��R&v̿�}g�1SSa�
+��~�;5�d�PgP���p���Y���G�q�M�!Fǳ���w��4v� �1HJ �4}��_9������7�s�=8�'����iv��Q���U)����e=>�}���!1�BY.�j���R+i��r����9���ho2J�Ф&�i&����-ʷ�Wv�~�Y����Q@HĦ�4�K�޾~�!�����Ə�],�Y�'T_�Y���7)H�m0�h?�H�:bn�r�p+?�.3��}y�6�g��&�a�4��k��H�،f߉x�a�9��04���F��|Y��6_%J�
"�Έɑ��c?e���r�4���%��6���i�v�_(�E>�}�4�B�9p`�(��~!V���5���7�Itg#��H^�5E�L7��{�Y5�˸xz���8��p�/E~Nd�o��,���� G� �8Iq��`D[X��ҝ�e�<C�����顁ø�I �-Tk�៻e���pbv��~0N��:�}žE�G+�}���C�S`�nfq�!�|Qe3n�â�����<�$y�=w<��)G���Z�(d�{� <�}�<�Nc�*{�w��ܮ�3<��Ft��Cݶ��і��g_��!�RC�}z��	F��f 2�+՞�����x&��w��b�D��O^n���I��Ƃ�OĻ�=��@I r�Q5�����/6R*��tI|
M�bM,�M��6|w��3'��q�N')��sk��Ҟ�hk=K-�-� ���pr�Xq��|�9oP�T�}�P���k2L�n�1��-`��q�Ixao[~���b��'	#_�=nP��2�
-�X-��QlTB��n90��p�"�K�őCՄW��.�/���%����]��Ӌhy���&/}]�Xw@�5d�x�=ף�!�2�qG�Rr	���b�pRR�v�d���<��Q��v�H!�U���]M8��6ܘ���M9
����֮԰^ ��/�E��ƥ��Eik@��+�^�+VhpVYD��]#ב�b9�\��ڿܙ~#��?����=���y�-���H��}�z.E]8���|�߰g���كu7�8y��-��?�? �˂��w��C#\߭5*�x>Q(ƶE����f�����*9��/�#�o�����6�����	�
�MVza��Ц�@���۪�B�Ts@"���W@0mj���z��?�����IS��$j�;���ܬo�I�Z3��<��ľ��-N���z;��%i_����fZ}��F]r��}�4	�|�`7�5uK,/���d7��a�I/�Xa�K��x��1s���Hѩ��	�\G=�K3��,K��c�ۣ��d��-�WFc�/"�0��(�sJ�}w0ӂ6�3��^sV(��*�`�!���cӠ��Wd�*�Rj�iuu�u� �/i(�2
�vFG�9r&��OiH9�Y޿v��
=�պL$�Sғ�I��w���V����J����.��*9�5�����"2�Ee�{�SJ��0ӆW�����9�@?E>���#\��u�>�cܭk�r��2�>Vn� q���.�K=�麢��3½���������@���Y(��m���BM�L�Әى��F�Ƿ2>}$�D��*TB�r2��N ��|�T���)ӂ��+z�]J���8y�h��Iǝ��ڿo���o��qJ�&F�Z��ս�>��9�$
�^�1ճ��W��5���E���: W�|�K8���5����#�<^<�XoHM!9�3�m��8�Йz2��T�#��؊e,7�_( ���N��a�9�]�9f��i[1!�| 	s�6]��`�#����'t��l;�e��������L��*Q�iRa!/�I�.��_0c����m�3�$�Z1	A�% �tR`�f^��f���G�Ө�L`��*fݻr�z�b>َ�����n�������Yx��p�[�1��[���4�]���:1s�L����0·Hk8l.n�6�U�t��C��2������%h̓��ޭ]d��Đ���U��r�j	�L.��O0�$l��[F�h��q��B]��x�kQs����3�|�H���P�_lxt�'m��,(���SM�*v�|k�?D��µ���7u��H	�B����ʓ�	Ra�^%x]<u.O��$���� @ul�Y��EFP0]�\"Ri�"O�Ռ�>�#��)?�^Ch�."���%���P�l
!-��`;��6��K���:`A�n���:�=Q�^�<�#�O]O�$���a����(r�L}�o�zK��o��0�2 ���ˤ���aY�<��]�!λ���j��^�O|�MW��&=��]hc1���@���x�#i)���)5��/�ܦr�P�9?ֲ�1z���о�N�$�lP�CB�ht��p��1g��1,әl�&��U&u���Z�h��k��P|Nv��N���$���˂��n����b �M|��ơ#����(����ST*.zؓ�����u����F^�̐Wx���������4.�=,PՇ'v�,V��b������p�I��o�p�Zj/w`��m\������᫵�����{�*C'�A@�Y�n<�앨��5&�w�
��E����&߲���JŬ݆�*�MT��T��Y��PE_���T��̌VS�	���]�]��Y6���C�!D�Rf0���55�9>�r��3@�VȀk�&;�&'f�o��j01ȋ��J|Q��9���A�8&����m��.:��}8 sL�0��Y壜'��d/Id����m�GW{{���Qc~)yI&���+�Zz�������dq_��hz�X�-����x�l�?��aR�����aQf�'j���r=s8<�������� f�rT;�#�e���>��S��gܧe���>�ʩ5W���z��`@�/]&��C�� W���[
������F�n%��eF'��9\�D
��ߞ\��ZӿF��QQߡ�������b�؎��tMȓ��0' P;czڑq��xI�9���}��Ή@�d@�uС��+�^��J��;=��r`�Np�T����?ն�)F��E�"Xby�k;E�7/hN�e�F����uU��V#܉�x�a�qh���m��7�J�rߟI��f�b���|B<ȤIT�k��n�� f)GfI�PM�ǈ�<�����v+���-M�
b	*!�y��UmX���|[�����*�z�ʧ���-�����9������$ ����i�1R{�>�.6��M�0���L4B�dZ�T�O��&BN?�@@
1�����
ޑ�U�_
00�m��0�9s��D����8 {J1K?"3�#m��<��2Q�F�Ќ��^ʻs-g'�X��^>�X×[��f����6�؈�c����0��ʅ�Ю���ee����j�*j�q��l��CJ:�d:�/��tj[! w2X�l���l�7P�����#	�u�@4	B��V�^�li 橷:�R�"��f�Aw�y����?����Mg˃��״9k:������f>[������Z���Dj��#�#�>�2��\�׍��D�Y�³U���� _���KN�(WsY�q������d���UX#4�.��6k�4{�$�m���Km"Y%��iA����.�|����~� q
l�-���2��з�x<}k_��X-^b%��ս��Of�i]����T{�͎��j
��6M� "��q�����Ud��N�+�LR����2�Z�"-a�]ŎgVo��N�lO=M'd��%?�4��K���BU.�>B���txZ+ ���w�T;����χ�}͞�� �8`�MoC�$Wb���Ez��,s�#ob��QP	���N�IR����"�%��D0��u����6���A�H=�w���r먿cךW���a�A�N:��sZ�	����w�,3�HZ��E�@[ib��#�K�)[	;5���՝��x������BcS��^��A�P�*<Q�kj2G�]����h��g	��7��6��қ ��d�*~O�We'�����O�����\Z��G�MԖ�1��hӧI@�dO�ŋP4ڇcԍZΐ�w�S�sWd�ܥ�Ѵ���awfhyK!,��@�#ŏDzW�4���f��v^Rn�=j�.:� ն�f��B�$��eѵ���m��B&w�4ሱ�䦸̿{$ê���F����l�6�Ci��!�
it:�[�̪��>��٨>��ܛ�z�?8bojg�T��\��T�-7f�������A!���"G|��(�&.O\5�L�8�n�fg�o_�1�����7t�(~�J�ɯ��~\v�!9/��}�V�s&isjB�	%Hi� ݝ��w�+�i�XS̃�0{�0]͒c���� ^n0��%�i�l��%Ugx����8\R̅��j s�zIF��ŏ�?E��º�3*{$��B�T����A�`����gf��sѠ>�
(�����M8n)�	��`L0A!�-�`MD�q����]�π�25�LԧL�byX
��.����7^�H�6�~[���{�_<=��pͺ��K7>'��n�p���B!�-t�5����vcnc����խ��Mu�#w�U��oMng쮉(����O3
y_���XdOD���5���Az�§F�Z���<����f�L|Mj"U�L�3+(c�7�zP�V%�CYph��-��.R4��,v��.�,�Zt&���r��yU^��$&��(WqkE���˺�l�?@pߛ�Ϳ�vZ�p�B���٠P��o4��sd��@Ѯ�f����ϋcn2�/2��9 ����kFږi`!�ƨ@X�FC��9̿�21~hO.e�y����Wzm{���I�ک��4(
r��o6���2�e=Hd�M��G�ڙQ-�\_�n�e�Y=����n]\Wf�צ��d�Tb1>����u�DH��8�6�®^am��kB�-J�	5����l�϶hȿ��ķ�ϣ�5r�DP���J$��w��D!��)b��%8LDS�fvUo���R�&�}U�]��c�1zJF��VW�^�>�]a�����u�X;) SHW�r]Z%J�R\y��Ҍ;��n�׋������@��V&��NU,3Q��<e��m�C����/���Q�5E�n�>lH�4`��G'D��ΰU~�)�BX�?%m��L`.nF�$P�^J�9V#��P��I^YI}�~�̐�Y�_�$��#��Ⱦ�@�Y���/pg�ԍ'?����v�q�R����N�{�T�8�U�����o�;�|�*[���n/�򰺾F(I_�d���J����O���r��w P��R>-��q�g�YDk,�������٫P8�h:�zͧ��i�|幦���¬o�Z���P"g���=�d�k�RW+e��U B�Q�B%a�w��������adn�&%�����#m���%�Dw�+��=
��j�h�A�yn4�d���[�'�?��O��[�w[��c���N�>)^��鿣�����x�C1��3��?�R� ؿ|���f�+����`'+���������"x�'��:�3���j�(�����y>x�mc���>[�ܜ+.� 1�s9㍠�N!%s�8{P|x���I��/��(T�keVE� J(n����2�N��D����Ʈ����6U���h�6��, &�$�t���ÏO�,����-Cg������B�QTo�\��f$�-.� �JD��{�y`�t%�x�zB�Km�/��>N�9E{���Ç��fA���6Hć
r�='��N{�殆��*	*��4�2��g��@�z��ւ���
�Z��ע5�V{���2�s(��H�������dI�lEf��� EA8���S�����#0`��I'�;E�\w�w����I�}&�<��]Vh[��B#Z#�a Z5Ӷ��i���x�O+Eq���޿:��">e��g�}�\�Z�\���ڊ�����P��X��3M$#����a�w��rj���9]�:��a�YBk�����C"�W
�����<z�f���)pOM+�����\�e?�`�m�P�q���ұX���!GX*��f�3�;s5�~�s��6�
���\z̶2h����K�6BC֠N!�6hB��2��b?� V�x�ۑ�����|�����m�#H�v�y�kT��H���$`x\��/*"<y�/%ao���|ˀ�vO5��ZU��FƖ��Qo�sQ�����Vr����E���.�6��m�x@"�(�ȗctn�6'D�����J�M�dzR>��潕����bU%
��ߒ�5��pq��C�Dl;����, �����/+ؕ�G2h����
ۤ���֎�1�%�|�����ԘM	��_�.^����̱� = 4ş&�D*�F+�Ԩ��`�=����B�v;q �D����&�@/���Q��t���\؈�@�ab��j闠����LU�rg����v'���"��A��P!��/�5i�ͺ����>�_�i܈��'ӓ;��<T�� u*%�����`�"��@#�\���腑�#^
CYX�����,Q)�X���9T���]MY)~Eо�_ Pm����/n�ѹ���Y�*ˠҌ�!%�q�!pX\M��22�^�ʱt\��6ma�w`�Ŝ�(z>dU`%'{�[�������S�@���h�*�~�rF�i"eK递ƑRaT:ˊe�^��$oz���!d���gĴu�q!`�s��*���AE�ƌ?��&Z>N��
Q��j�+�:��aw7���|�-�T�N��ȵoN�3~��O3�S��T=p@��@u��G�eE9�k+丌�68!�9��?�>l<~�Ğ�!�ٓ��Yz0w͒��	|���6�2f6�)�q�.�����Rz��,Ml�>d�(;�N��B�j�ˌ��Uq�)h�<��nR�7P6 ؊�4.IE���s��.���?{��z@%J,+�؀��0��czo�(.�@ަ�N,���4m���Hqo~ͤ���d�iV74<!&�vv`��s
:��d�����?'�q���Ws��s��	-t�KjV?.5*���v�����;kD8�p�aXv�����g��ĞJ��@p�ԓ��/��>�J�X+{#���G�>����:�������sƃv&�Nm9/�c��g�X'�e����o+i�r#w=��7R���@(V�o�;#���Y�J�S��ex%y?���z1tE	hv��Cr�1��O��jaw�w���"�TJ�\CA���@B�~G:��a�@��i7��e�18��	p��<-��e�I�ҵFh^�ty"}�]���=�@`Z�U,�bh�y6�D��p�g�^��|BspRF�8Ako�`H�2���О�J�,��0����->Q���wJ�|��#3ɰ�q�J1��<!�=�k�a���@�b��O�ņ���NCc�#����!Y���([�W�%M�l�G���&��(�Z?V�,Q-�ᵡ�|����W�~�N��Y*N�F��`,�ؐwi��A�(N�����\��nE�z��4w�ZU�`�f��{� ������Ox�ۨ�m���!H*���=���z��V�>?IF7��4De�9�έjR~�̺����P�]N~��1C�4�^sS��\�Wg�����mɽ��2�2���fhU5���}���K�,�N�Ycm�^ա00�AI~k{��z�R:Z���L�RՔ7v�}��أu��g8����0z9~�V���@��/88��]=C�WF��}� z�(G<����=R�#�q=)xgN�9��.�Xv:yd����MN�hgS�i^p̋l�6-�I��y�Y��ы˖�ӹ�@$�nl��8�ҷ��`��Co�`9����r�͚��؜�����#9e�I�-p��6�����'.���]�K�����Ù�0�묑�,����oY�꺡āV^,�'	���	W�MN���٭�����5�Yt(��u�=��q�4��NR���,x�/5���X6�5x^2n�wչ~E�Lz`\\��s�wN�c�i�*#�la�ے������{Ab~I�zdѺXz��-�O�������"�c���������M"�mR1ʈCc߁_8 �B0b^��r49��F����IW=9/����y �����Z ��6�&�e��ƒl� Ȯ&�<�2A�uP7���XvWg �s�6Yps�/MxRd�e`��Eַ�k�P�b,�N��U�h�/�ŗ�ˠ�v�-yXF�!�I�/�?-�醓+z}[�A����MS��b�;3N�[�O�h������;T��kI�8噵�� �
�����Q��gUM�Y��[8:U�c��<X7�k���F��Yr� J�.�澦�������a�},^�Xn��j�w"�O ��K�K�|du��}%�����II��o#~
w4�P@1�%=C���1�E�)�g�&�6� ��{ ߥ��n�.�Q���zɔ�ϯR�n���AӇ�[����FS~�Xr*{�J��۠��%(	�㙋�=�5��.���Ƭ~�%K��]-�E[���vș���8=|U �,��m?�.���Z^�Ր&9U;���*�&(��������K�?7�kA4W!�4B�B]=g,P�R��Rs���1�K	4(!�l����Աl�~K&��u�/�N.� _�:��Nƭ������0���7�G:&�T���VD��u��{R~ق)6c�n�&%v"Q����t��.���p���{�}��y!�+��!y�)*�����i�N��7{�dd�7�/۝�;���f|�]��ɦ��n��/��*JH)��Sg�X[��h������1WƎx�F.c��荒�4w**�Q1��%HL$�w�c~-�Yb�J5dE����7�˽MkZ�
.0�Ѕ���TP��A���<]�]����ʝ��7������6������{E����o,+�)4�͎�b5��%}}q^�l��
������l�b���֔��&~ i��q,�J����}2��ɦJA���AH=�����Ǖ����X;����������h�q�{SwyK�.]��B�����g`V��T�|��V�n�/u����ŴS�l�m��\�c���I[�����Œ-��@�|�P��Y2�U�(���Ф��u�p��JP����D~�CO)�@V��I��"]���k�E��'�&dY��Z��ro�(�8�a��pE;7���;�C��L~a�@*�煯VS������;� �D�w~�C�\��$`�
CG��aY�6�^'��s}�қ�jتeȐ�W���=�^F/��<h"�MS�붑X��) � �F6�ҿ\ۃ�x�)�B���1�����@�̼���%�
I�C�2A�<��IIܠ��x�:Z�(����~]˫e˪��~�/Lv~V)dk]T�	��9��_X�"!�M>�%=���rɘb�A.H�t�+y�# ��<(�H�$Ct���R�:@/��N�N%�&J���`P�f�b�:�J�0j�W��P	{B�V�Oi���ǰ�9�:o��4w�����=�-���2)��0���gTcs_���57�61�u��������TB�*Y�x�{�@��KT�Sި��#0Gi�9�Pp#�"��(�t�+}�*�^��ǿ��U����dyO��Օ
�͇����Fj�h74�Kv��q��/�i^��O��2Q���N���Ω� (Y��V`�B�����N�	6���@h���l){���u监z��N�YM2݋t&�ޚ�.~t&�ŷ5x̌�Nr�S���i
HVT�r${����7��\vb0�^R�������;��W3�!�ًKf��Y��-��"�x=�-*D�f�mHڠ7,3��5�5?�Z-��+���*��V�@�M����
N��Q��2Nt�Qqi�'��P:��pX#�FO)5j� '��6�0���N�����Zw$���u��X*���������bB<zWR��γq��=�N�Y��0��w�����'WA3�������-+U��jK䌰
(D���R*�d��1��n:XaF!���+�$�X^�c�_Q�V>��3f}~�>����U���eKU�[��>m����;c�Cʜx�-�'$y��}NM4���敐w�ᘓx��c��&����;�p���yO�u	��&r�wA
X̩��W�	8����(߰�x�B�J� ��1&�c�����ѭ `�Ҭjߩ1~c⮦O9]Q=j�f��'�nF�}�b`k���K�����f<^=�A3�I/���X�jA���v�HS���In��e`�U}�o#����/��b�a���Ƚ�(�^���ތu��K"��)iF�Y�������}��F���-�.7�?�=t���$X^�����Z��讄OH���ɡ.Pv;&�GWS����*[��V�,�Mz�Lc�r��Y*O�_���9�"�JW��*4���|�|��L��Da:������&�:[�g(8X���#M�;��������������ܟJ��Ƞ��p���^����|D\���B]��\�>}�R�i%k=+(��ų/�!Z)ꋾh�yQ(@��"�DD�Hs#膠~����\A��8���T�51�/%?p�� ��H��;:Tn���������ṅ�y��H�&0��7��]� ��i�����)��C<7�fd��E�C(Yo�Ԗ�C2�K�5�JQP��f�`�%q�*�N�dP>6�@�}���(_EQm�Go�J6f��/t�/]rSל����w�?m����UʕɳTsG�p���**>Z��[�ӏAF 8�,d;ߪG��A� F�%�k�Ks;-�#� v�eܶ@���'n��qV�CRxv���%��|��J���xcm�+��t2�G�.�^f� ���	a͞�@��+��H�yo�Ӥ�C+�<OB׀	�G`ZF	�Q��`*�,��X�^j�$nx4�M��� $�d�cµ7���+"�|:
�7���o�dLs��N!>���*	�Y�z?˦��'��l]m^��_�ZP��D��\~����A`��ZA���K{>�=bZ�Z��ļv�(����J|�V�����~��8��[�Ēe�Sg���L��m@�~��f�_*z���(�ls�~�K#U�����ro_��uK3��x@%A�2��kZ~����ѡ7�
�qj���������X�va��@��P��o�M�#w��Z�im�	vs=����������X#�hz��q@�T!t�tj��?�IUc��)� āD�rG͒����?͜�a(=�I4~���;w�>B�/p^ckpZ�M56�v��A%[N=�PUN+����b&�Xщ>��"�h���y���lԺ�����1�N�8@-�� �-�=�[�=.�V�>ZS_XV܎T�:�'��@�OL0�k�`wY�-��b��{jE�\��������/v�n��x9��Q���/u5��o��]��%�76�q��_H�q�	��O��
�C�q���ك{G�<��>�qR�,��K�Z�t�CQ�"�L����S)������{[��^�Ɍ���N�V�-�����~&h��a�_t�B�Ҭ"���ڻ�%�`I�Q�v%�6�o_�F�;��E�l��k���a�9�$|��I=�Q�o�`5P�G�p`.���f׿m@�A�e
��$�B��C��&���Ew�%Yð�@��6����V������d�Qt�u����w�2���1E9у��I�f��~Rc$�F�r�`݂Z�����ȢC��
d�̩�ړ�܍S����`��%��#��vL�`�B��
X(�j��.6�a��l����2�;F�m�N�j^d��m2ئz��c�5�¦�M����[�0��6�Cʝ1��?1h9��A�3�0 U|�Z0�RT�!0`Ӈ6�X�p����Lg
�����h�L �;��n�QMv�$m9W�sb�P�
c>�S����l�t,�,�-��ByZ�z��Y�;�⬚p@PU<��p��=:,�T[c�sU�!1�W*5"ؔ���&&��?����F���T2_T�<r����u
QO�0>B�7,�ngW�%B���ǜ�$	�&L����-��$(N�/���.G�]���t&<?;�t|G�k�PɫK�m�8ۓ�SfϗC�x��'����Y��EK��&�!v�o�{3��,R���c0�0E���̅tсpԧ��
O����`/xG���S`����T���bkS��b$�\�s-C'>_즂�cF	�6�DO��Vm'մ�u&�\���NW�N��Jz�ܖr��1����r�]��@�=��a<��|�7J�<CT೯wVk���oaW߭�)C>N/��Dq����<d���|4_�U�{nc�#�(��q����x�jxt��x2�:
1�T�^��i�Z�5�.��֟�O�������	}!mv�O<�#����-Y�Q��8�b��t$Ctk��6�	|��>S��}���,�Z?�!E�F�7�1Ѻ"���I@��fo���F\,�&��ysU�����R;A�f7ގ�9u�a�^�����%5�dr��D�em����~�� �<����,��J�(d5#����J3�0o-
3^�Ƽ:�&"[F�i��.z�i�Z�L
�u[n��)��U��|H̤"9��F�[! X�q�-���Y�a�,DN�"GP>V���tfPM���j����p�
���lmE��E��Z�D<��I� b�+eY�20��92��<[{��^�e�t�=��F��y���d����2�w��'���mU�q���i�kYew���27�M��;�%�,'UN�-DB������'�Șx��ToD2�iݹ����-��'����lm| ֵ�眮&�r؛�� �ɚ0Oۍ��RA���Y����Q"�mM\�=̌MVaT}t��DXV�'�����|u�"����W��t!����'��F�UH��΍W�>�Cj�	�H�V�Y^=V"m�'y��_�`��͑��r�g��6@��?)=�7����u|�����GXD���>��<:�aL�>��u�]�M�MEY/X꣟���=��,��q���[#�Q�HD�"P�f�'�o'���-���_Ud�+YX�#���i�Q^?�X[�>��>�U��W[U�8Ì+*H�}�[n���,q�RxGB�2#�hh�~�n^���O�B�ۀ��ku"���,GJx��"��v�N�ګ�Ƈ�3P�%L�Y>%-�g�t��$�~%g=�;��1��G0wzH��5��5Z��I�4�!H�9I/����S ^� ��"Kf.�<_$+�ʱ4�F	�FO`o�)Lr�Žy�Z�.91�Q�?�w�� �"��15:�)$^vI������~��*��C��Tn�����FAY%�hw���-G���`*h�l�@��in S��\͢�D ,,�`��R�ګ0ֽ�e�A,��� 7��6CE﬛	d�H��aѷ�F��I*gJ׃^-�٘����ӗ+�`h�/���:��~�����W�qԭ	�Z,O�۵m�rZeU�'�w��P3^r�S �x"S-�)�h���q2��� �o�]��5X�Ki\�}���6�(Ko"#�,I�h�/D��Fa�~&�P�8��/,GC���ކ��+��h���˨��u*�z�V ,�A�N�c�}%������X�;�@��9j|z#�N������7��O40S� �6�t���b7ﾛ��u���|o�~x?�̋$c�J����c%��SW�;v�a`�}���P?>^u���S�g~�;�dS-��"���(��|F��}ǇG�Z��{��#�ݟ�BΓ)}DZ,�۹sYy��30<¦7Y�wb|�}�2lB�(�Q�S����>7�|��tR�%=S��.��O�1�؄Ji�Ao�kvϵhe�ˊi�/�@�TXbAv�v�3fhJ���f�Z;T�Fh�2�{ݙ���}�K_�����x�΁Z�AIaS+LL���e^g��剃)k�����"�m������FJ�"�Kש6�B|���{S.�P�t��5�v����,��N��%�-' �&�ڶ�,<�G85r=N���Z3�����~�h�'�V{�:�>�O���vڱ~���9�l�:�K΄@ˤy� S��R ��K�����xz�:N@����'��
���� ���m^�6g�z��LJ �<R����C�<'4B�Y��%�|�WV	���2�m�h��YL!��1̶y�HU��BW}�R.���d
�ut'QCY�g�_��e�T;z"�s����+tsK��$5_�l8aj�*�A�
)�(�j����
�{vj�xgŀ�޼@�Y�۷�<S�3�n͆wMmm��s�k�Y��X2"�μ&�;�#@yݝ��e��5�)R�5
�d�����^����;�3���v%����^�8��ub:A���ԏ+б�2�\��Q����1��$DN�~)���5�M^�b�-���⅔S����U�M�a�$�=�	���B���?Nu�q�S���Zo�F*�Y*�-c��j�g/�r�=(�e�|��3�p�
�
?�k�ܲá�6_��rی�$il���N�w�⢪���<��E[�9�@��p��+T�E����oJ����>o�L��;J��dj<K ;�A���x���fo8U$���x� ��&����oA?^/�O�G�=-��	u#��9�R����Ny��+��f:\���6t�E��3!T��V@&�<.�;���en��o�mT���F5t�"�t�YF4^��T�ݘ+U�}�������ԆK�p�\��q�E6KQ��,�i�_�[rΐ�~&�̼q"`�L�RZϊ�b>+_��V����<�?��/j�Z�X��q��W�l�1�}�b���S6=�V�n��כ�i��h�A��ծg�ؚ�.nuHE}ƻ�~BJM�9�(a�k�{�x2[z��!�ԋt��#v��>���n��T��S�4sU?�֧1(G�!|xL�i%��l^�҉�Ã�l|"�c�p��g�F�*5-�u+�mY��h��J�T���ټƛܛW��?��F=э\p������vE�ge���7����jE�a������g��iݹ����� �����1��>�Q#���b��%F�=�s-E���e�����U�.���$�,]�.�/��Ȁ[���ϫ/���*�1��NT�<ʤ*�'c�$�� �p���15n������8���E��c5D�XL���ᮩR
�R��۶�q�����X����_���w ii��hz�!vL����]�s7^H���L���9ou�L�ܷ]�X$ ��ձK�%� ��q�o��R�Z���%1J�Z�&k�P�OMf:1���X
T`�s�ј��i��4�2� � U��%z�c
�����=���=��TWd�x�ں��p�â�!	pSW_�=,!7x�e:���E�2���	`�1�nG۩�����M�
�K�cW*��y�"�МaC�%N����Ub�B	QH8w��mFK����6��M���h�f|t� ���Ar��<1"������P�����.<MA@�����֖
�D��x%����F�|��F�m�"��U�AO�|^cu�y���&<�L�"��@�
H���\	Q�����b+}� �t�\{�t§�/��N��I8׌��߅�h���S^M����e�G�(�=|��.��V>��Lp�9r�� �՘]������j�G̸,��~<6�(�]���+͕�h�W,1S��S�X�_�<�.�hm��o|�QX��r����N,7"z���#\����;H L.z�	����n����t唷��j_Z�9�A/)�S����+�Z�#���||$�j�R�XnC�u�!����}�U��@_� ��.
ۣ�dk0���4e�o0�nax���Nc�|ӨF����t,qo;_�vm���?�Xk4����S F "�0�њ�zq�&u?�:h�)R(���;V�k��@c�.76 ��~?�~������1>�!�ĺ���"�Q�_���Mqڋ0�i�{ȕ�f}���4ZD�+'-j6����z�i��l��L��c������~T^(�W��e����<�= /�J��?K�� b(<Jn�������B��~�����=���8��ج5w/�!��d����bv�ɏ_+�Bڗ��U���i�;-�úX�χ�#��Կ$۞Y�܆0���B���TY"� ��^^�����N=���B����w|e
�������b��G�*�JLw���SU�"/y]k���/�����ڧ�S2�qS�i�u��<����km\'��&W�?�4�`u"�[Q���q���dO�T��F���J7��b���(���t;���S�J��{���M�:���p�I$5���\	տ|�B(�mz+��YA�D1�0
S1p�L�r'@L���P��Tvџ��B[��`@Ad+k΄�OG�8M�7���S�f�bIX�o{)&�(DL�R
��l��0�B��RS���7��>�Ϝ�(��sӔ�)R����7oq�J��O���a�z��N��-ͬ�����}���s�{.� ���"I�5�.v��F�����Zi̖��q�;y�A�8��u���������L�}�%|�@(�$L˹v��B ��	H�`�2ދ�"���3G����N~�	!��zڋr>E�����Oft�����V|W�!�	���l��tt*<F��z×%�9��/�Φd$�� �ܐ�v�zMI��ܻ�%ɢ�s��wl׶L%k��ꢞO����sڵ����C���3�]����lQ�x6u�G�u����Y�~}�o��ޏX B����|)V�`�����u�x��Wt_P4�#��q�dHC�L����#�aB��S���l��!��)_�ؘn�_i"ڜ��$D�̝����0��3Sv�@0��x� ��wd���������-@�II(b,8xߵ������!�5v�G%J�Jǧ�!�H��fI����d�l+t1�����ܻ���hxE=�������� �ʏA��.CQ�|q�\�� ��fIg�R�İ l3��鑅=��$�t(wI� ?~[#[�;���M_�%�_-���, Y��*&Mi�:VS`.�H��E^@�%���Y����W�h5a�`P�\��]q�VQ�Ab�]@�*.�%[�K��[�]F'�����v���s�;��Hn	�=R�"���v����C�*�{j�5�)�`�gۓ.J.C����y4[l�`� ^\M@�����L����!c�&�I��N[���>׈!4x��,���HY�gB�#>�)��%�`4� J��kE=���40�~!e�"����Nd�9����I3���7�RQ7k�π�����i}#��#.I�ឲP�hյ��x�iC���&6�x(��" ��tlqII A�d�A�� >���į5�7q'g0�+8C�
�8Ԕ�#�����R��sPV_�L���%���R�m"���o��Ɔ�c9sH{���? >s�P����:�teI$)b\P1��_r̣r�HNr���F�#l�u��6tn&���5�n�AӉ�`9�x���[-y��y�^wwqy��ً���I�E��������m��	#J���S�!Wv���3r�W�R2�1��wzL�&��G! �등���`��㉗�m��7�x�LrsD���m�4�@�2� ��S����_8ڥ1��Lk6�R��t`G�P�6���A�,��1��Fصy|�90"�ݶD���\[W�#�2�I�ΝV�0>r��i�ov���_m|9��O�ŏi=h �-/��a�Pp�iX�U6UX�l�'�MX��]U�����yM���� 0�x�C�i\P�5�sc^Mg#ڙmMLf-��X�x��D��#�������7+W�)��R����h��V pk��}׫��)ZLH�i�	|��%�Y�q�D�+,x��`A*@�_jf)<��^���,�j�ї�i72W���v��Y���.r%w�?�r���In�r�->���.?��� ث���]3ը�4Z����vy]��R�3�:����q�;뾼�T��U�'�V83Z��-k�IC���].;�p�����E�jr�o���1 �w�����<������QÊV�����u���we}�����8���T��9c/Y?>�o�����MT�	*,:W�L���������B���+�}���-�2�s�2glv�q��c�\�A�.L��*�1�M	�;�DgDM�� ��ޜ�Z���(�}U!W���"���y����+~�MqW(>��>�&M���$b>b���Λ����B�y��b�/�h���A#WC�	�?�M[�S���A����9��1\Q�7��l"T��6���#K���AF�⎃5���?D��`�qB��D#���ʘf~~�T���G���{|I�?Zt9o=K�n���kԡ�'��K~+w�|m���|�&�E�t)�XVe�;����xr([�i&��s��.P��{#��WR܋8�HD�/r�<�淣���ꌟ��&q����`
�1�:��z���$2���T�	.���X��?�6�/07�
l�P�2�/{���i��كe�e��qѼ���B�u�?cWa�o��M%IMʹ�v�~g�"�u*a�{pC�?�)x�e�<�|���@�c���.l���t�r�e�Ⰻ�u.Z�5m��ab�� {b[}�� w�JW�A��%f��pjX���'t :�q�<Ѻ�8��"P<�n�XZ�v>[���<��� ۀ˪Lʉ�_]4G,�3Gx>A���^�>m !*���_���!',#�&��U��:���n��"ϙg��R�*�p�nv�|�Z�K�41�_���&!����܂i��b�c��풰2�睙��_�i�� �4C��Zkb��ۏ�1�t�X��9{^+�i?�^*��m���1���>��B�C56-� _��?慥�5 �����p�z����`��Z~��'�Wn�	fw?J�~�)ܛ����"
�#Comz��O�-���v8o8zsB�!3r����p��#?ѝ��iE'���R!��K��>; �_�M�C��?cq�=���~F>'&�h���4xzY7$̰`��/�c8��i�'��4��]� ��=tF���s�P� ����򔇜���PE�ܗA�a�����|j��._�d��e��h��Vf���o{�(3����!���P�SE�$$��g(�T��b��$��V��<[j�7Vf�/A��(@��?���NNv,���;����\�y㌵6�$D���p��(��������)�3s�?�_�9��ߏ��B�.D�>�ά�9��߽S32��!�>��s9�t�Le\ݓukC�X@�wO��&���}�+��₢��zbM,6��{���R'�� ��
vࡗ5�v́���3��Rl���ڍ�V+C����E��sީ��W�v���}�#��(�%�Vڶ��:ހ�O�2d1�P�jNP�ciO\��_�Ӗ�$T2p!3� ����RT�Þ,{+��N%�_�_;9�(����u���<�Jۻ;��"M�jH'����"��h�hL��<{4dD�*'�I)�@�Hϕ��g�JZ�r�ݭʃ�����ULe���@U�Ӄr�� W�m#[?�Q����P%��Q�����z�����\g�_�j��#�Ы3_�C�A�A@��jO%>�t����Ѿ�!F�Bg�?Z�k�3��f$xV2��ST�rl~r�����j`���y���>�v�9�`���@b��9��i$�]�a�0�&����*"ȤPH��� ��?�VL�ԝso#�� ����S�Z�=?�8OJ.Z�CF�RO8�<
py��d�+γ��Pߡ���-��"�fg����~�!����H�*�6ՒHI�r��z������wM'��5��7y����x����OY�#I�t�2\��c!���f뺉u�q#0Eu������l�p��]�N�S��_A) �x��?���>+�\�(�l���M`o������?!��ʯ���A$Ÿ����9e~���o1�z3n��2����x�:��̀-��ܭ+�?�N�^c7 ���A��xr3��m�ž�G��$�v��0��7{�lH.����|�	u��SC-Ӵ2��(j�*���
׏rtJ��>}Pc�S���^H)m�2|����������I�*at�Dy#�6`l�{�5�/-�$ty��AG��5}{_A��Ġ���/��a�l� ��9�G��}�!+.U�EC���a�57���f�AEF���8So��to��߯7����H/���[jA���: �
�%�{�t�M!���z1bE�m�m��9�p�	V;n��v3���@�����Đ����Z1��
��1���J�d�4cf|����P͢��#eWCM?��nC��QG�Us���Z&���8�?�t��k��$�3Dr�h��U���j��m�a����3Ǆr�"��f�>�+{��Ŀ�\8X.�qFҝ�25w���)z�Kp�DS�l�EѶ��ų��щh�+_��]m8�h��d��|h7�N��r�qS��8�k 423�0ӹ�
Ԩ	2��'�˧ʲI3y��h\Cb}��~�ŏd� I�7�f~��3П�Z��N� L#!��*�>�|e�u�C���.c?m��@�H�|иN�t�����e� i}���n�D���=B(�������u:w��oq�N�
�Z�
��xǱ6B�E���_�z(	]�0"�Pc�{8 �]0U�0����2�p3f��OU3��������iEj>���V�-��P�?��X�nL�7�oj��O�qQ�6R'���F��.%5u���V�
\�Oɔϋ�A᫂
��&�:Y�}�+��.�$�'�-�S�R�r�
t�U�;Tk$׎��4���c�v���ܧr��!�}��X��b���Ӊ0mmv�$¶����8��u/�����E�ħX(�F@qG!Z$c�A�c�)����=����re�*��$Z����K��(���է0����>[n���[m��i"������vcKƒ�{���?�Ř�T@F���yG����0pW>(�Yl�a��(s����˫J��^x�l��%P��w�.��چ��֌��Un�~�f�_=����!��Ķj��	oվ*4����(���ǣ��ʎm����M�@�f�Qa�,#���hϔ��d>�	�|�VYJ���۽�fA��_�I
MЫ`#2�Lǿ9י�%�����I���Yp�i8K���O�]j��1dB|{���tl�o�� 7����/d<RPyr{�>1�����Ԅ-1/�1IƌʈN�Űƶ�"��Wy���ډ3K:5�4�B��dI#�,n���x�A�5���vwv�,I/a��D�詼�F�DI�k���T+9��}=�.D��t��3�^.��X��>���O�M���{Y���1�Z�m5|��Ʈj|��1tm�v�˩��w��, #��3�l��B��b���K�����~�X�o�%1�5t��+�>q�#��7n�f���.B\-��UIj�^4:UQ��E��gП<�f���W6��!i ��kc�Sp4wqjN[9��	��7����;�O�f0�������9��.:�br���iR�I���lN��4��˿�;��K�;�ޗ��)�	���}@�B|��}jwAe6�؀ZB�{}�0$���w�0���s=7�Vh�`��1r� �87I&�s�H�R���]a�z�l�:����V�~t���	ҕ�T>G��r�u�7e������J�m)~es���ر>D�A��g]����$�6�ԩv�5���O]`6V-�e�@w5K|�5��&��C����?ȅ�L�[�]H���U�/M�m�'����F({_2[�cu�5R��&6� RJ���Kq�������$��q�]�/��Vn���NN%���: �;JCÍ�߬���0��w���X������>*�KX�������Q�m�!jk_r���!d	ŉ�6���.v����S�}��	&ǉK7o��댙�YvT��L�m8��%�T�-�I�È]؝�q��r�_"�;�2ZQ���S�e�9���(Ν�r����f��y{{4�G�-t;:�B%��R)�\wp��i��ɘ�s^.]����z���S�v��3L��6&a�#3H�����jA���(tA���O-�P�G�����<j��v�8����F�~U��|��t����?vx6��fG@A�V�W�n�僼��>�{��O������X��B�ə�>9\N��7�A���8� ��S��D�����gdKaꯧie�@)%S���X�8 ���y�=���	�J?�r�Yܛ��T�,�M��P�R�X��Of6����tY��'5�W��p�ȹ�qEj���Xؓs:��!h�;�-ܶ�6�D�����W�%7�2~w��a˺��4.԰�\s�1�����h����Eٻ4G���^ `�����D��i��#�߭����:$tش
5
Hݯ�4�M4����kji�*�61�����94F����"$Es�fl
(�iW	exX��c@b0X�������v����wӔ���eɹ6�[�#Z���^է5�9՛�m���*rI���0\R�EhH!�N��-(���Km3`:���/w`4�(�q�pt��8�ݼ�-�O�%�=��������d���%oA�I4��=�=l<����W}�=b��) 