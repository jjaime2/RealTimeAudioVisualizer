��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� ��5C����x}0���l�{��� �"�Du����!͆[��vgl��[B��2}	q6D�v����&P3n�hO��c`��`&�+&y��#KK��+�� �����%ϔ�)4�$�q]� 6�7����tLU�d�Z�����?h��d�RG�\��2p38�MLN%Z���1����tm�2�&�f��}����i��1@�g�����)��lh`��ڠ��F�=M<`f�r�Egq'�#ۡg�����X�(��Ԏ�[F���>�sZSM�\����M�)��3|+�� *x=0~���|��a��j	ź��X1�}mt����߇J(���j��q�}�@�Sq!Yp��i";����a\ޢiP8��{zׇ#@9�k�"D��oC)7��3�iH�>q0A�I��"�d��;����,z_Ӿ��4���PY_<�W����"G����	0�y�v���y��������q��z#�N��/��R�R��:�.��bZ�/�WA��V��,D��7�ԌR[tg*�H=1͇�"�"hL]#�Dx�;����"���+>�j{E "��u�E�B��A�)-��`-F�3h}'C1)��bȄ+}�9<�� &���H�3���nH�s�H�͌7I���~�,:����.@��N�?\��*8r+�񽩤;N)�,*e�-+�j5�WoA�P�ؿ��3�����G�	GF��@�z�pxI���e���v_ÔJY��Y!��IOt�2��g���F���PYT�0ͽ�����W4�'G�ꄇX����(�E�>�"�2�pjd��/��DZKo�6��.��E����u���a��(�OX��*�IX&&h���]T3{�̺	�����+й;��~<��V%�zU}�n��+�[ݶRޮ��?�'g;��#�mlW@y���y�
����^�7WG��_�v��~+��I���u�Q�㣍�-���KO��"��j^�o����5�����D�!L��D��W4?j!<�2]��9��Y�ig�ܦ��͟�|��.`wF�0�͆�?�ob�_^����H撫��MV%�)�u9=G�j�r���cj��W$ɷv"߸����M���Rp~�qz���V�t��m�G �k>Gδ�A������q6�)�w�蛤B�8i#JL/>Uw_�1'Rk)���4G���}JBX,��W��`[�vx�%\
&�S5��=����b3�QY�.W�$��sE�6VA;�}����i@4�?!(�e��[IU٫��|�����N�뎜�l�Z~d�']��#w�q�P�Ab��ݣr���}nyW$	�'f��y�1-@*�e���h���� ��i����i3��%�M/��%-���S�m�D�{��P��`�z��.�.�.d	��C_H���mY���Xa�DD��ɚ[,8�;0F*!��1 �� a��%��{�N	�:Q�K�/������\��PB(5d��\�����h����0	�d�d���s���A� (~gX�B\��������X��/KN�hF!]�18v3�k�C&f�$��!ӿ_P>���eƹ���^a�`�v< �Q,�@rU�Pc�Á�<�k�^Pώ�x���ð����L�P_�f�w������tz����o=��ko+#�EK|E��C	G�gE%���SƏD�2Ɍ�p�@�I���^�Ut�)������F`�]���IФ�H��o%�����~\����P�`��t�\���3Q��`�_Z`J*xaP� $G �A���v��HRܭ�����������`P&�"������@W
�oǄ��U'���������/=����ZO�
��cJ�oB�/��v]�T@��b9[�5p��RIV4:��ڟ��3x�o�IT�4ї�K�[ÕxXn!���\v "��1�ᵉ��a1�f�e8������ΫXkڻq��~�Z�(�����K	�4~1���ߒ�-�=D��|�ͺ~x<��X}l�W�<F+�k��2ָ��IL�6@��	�G[���D���G�W~y�g%a��g/8���\���J�OD[|<�h��z�(��l���um�8p��zK{�}�Ԍ$]�e�-��Md��dx�1=�K���{������ �9�{҂�_+`4%�[�"q|� ����aM�����f�F��A/N��@�'��xA^�r�9}��u��Q��G^�8�ǜg��la�V1����%^۬��ً�ɳ����$/c1����`Pe���d�WHg����Ô���B�1h��ni��eמ��v!�ÜE������00��NX������M'�{�!�1?�,��Vr���S��!��)թ1*K�6f'u��ÛY��SP׉���B�͝�٠hb�]^�1X~>�Y<��U��% E��!���f^��ra.�l�����9�OI}}ij�@�9�!u�NV�~����aeA}?]gι�/�g����j���|�y�߂7�˯��M�b`�E�jA�B�$��s��ijhg��	�m^�<	w)���b&Qj�>z}g����g��㍮>��hf�oe���5n Xe� �db�)�W��{eHޜ�ToxUJ:� B~�뒞�Zv�k��:˫j�1����t'��[�b���)r�(�BY\~���I�4X|"u�`�%B�4���v̵�	�ۥ�p�P��߂�'J֡�:��W� B]t9�U��i��IX�ӛɬM�0�k��u����'\���d�%9R��2�lOO�S8��1�+�}Ӥ���ުL�:c#�]0�2@5q��f��6aaƢ�w����&0�6����y޲� U1���D-��q�� &�Qa�+��z�;W�w�r���n�?�]�e��*�`��B����4����<�SD��L�70�n۰@�{����6��| ��Jҽ��D��5?���#%KiI$R�9�ޫs��57��pV�萤!V�ozK�7	������!�ez�_�̰.�T���9L��4t�	ʨ��Atz�ե�����g�o�8��"���<8@�� #:�u'ԍ�<J��3��m'`(̢�}���/�ry����t���gz�K�!>��H}��9H���je��ٶVО�1G����+"'�9�[�Wr�\d5���fv:=ڡ̻2r	�MA�S�x�d!B��O�E�Q�O���즎$ؤ�شN�Sy��2�_yV���G�M�#˜M�(o�W+���>GFT�Y����'���{���ߓ+��j,	YցO�^��7���V�C��J!\�lBU7V���]O��%�E�'.�z�Wc�V����\P��!@�N�EiOi���R�^(�C%
Yq��*|nu��)��7��5U�!Π$�.�I��Y`����X'�3>�@Ec��Y�FV؋�����a�ǔ�d3̢N��f2g���Zo6��-�9��4[��@&.C��?1��U�B��ϗ3���"�]܂���X�����\��T<����oot[�g�w�n�ܝ&S!=����5es�?OA����E��� ;���=��ij��ցp[�����(�;�F�j�r�*I���o���~��!�+�Y��L���2�����Ĳ�Ҙ����Ꮲ�^���c/n�PSr:G���
��P�HơNϮ����Q�V�,e"�2t��kq��p�y����
J6��(�U����Nj���W�����rD>hl��_L�m�:�'�������%�`�n�>�H���BD��鞇�NU@�4�/:4���AeMͰ�X/r����`9MX�Hғ�$�5�-ȹ�;9�-2턓�'�� L��vt�TԦ��@ɫ������Q���B��$����8Eƴ5]泷�X�FD�~�����PP�6h�n_���^�&'��ԧ���T���`����8��W���VFG�D�!�W�\z�W��A��N������*Qg=;��-�1䙾��u�+##v�}�`XAPx���B8�iE^1[	C��vT3��^c�����"W��榋-��z|�	���q�n� ����]���p�:��Yˏ���U�s+I����xzdt��Wy��tz]O�X�ί��_����q�cY����4�]�d�_��k�p�%�=���R���y���SlX��jD�$ŔH�H�(f����Gک�B��=�S�/��^�������t�@�$O��r�Ы��B边f $��t�"��Oı��؄��H�O-Wc� �Y|S���V��@�y��.��H�$��T���܃P�����͞�:��,"�R��s&�#�ݪ Ʋ��q=Mܿk5s��ĺ��������"x�'�g�?s��@�I��%i����q� �?M�6�
���妭}e>ӳ��F��􈚕���黦�|Q�]T>�ݠ�:&>�9�4��ӵ����-Y��"j>_�X<Y���ve�^���㱦�k���Ǫ��A�x�"�o��3v>(�6Hma�g�z��/V������6��+H�����׏����M5��h�v7i91&��-�*�wHj����&�"
j�J��T�"�8�hh� ���	Z}XӢ����K�@f���:.���[�ퟟ�5N�F��}NW�J�����a���U歳�9����N�hxX���}]�AbI<���3�l	�ā2//[s����r��ٷ�]���{��#lcv���oъY��;�c�d�⪈����	�E���ʻ5�@��-�3b��ZPk�d#��j8s��
��~��;"�Y�I@=���o,�m}i�q^�L�|G�!L�M�KH�q��'�u��"<��!\�Fq7�f�3��?�J<zV�38 �:�J�g�퀤s�������̢��I������Fc�,��)�i߾�U���$U��@K,~���nȑ	;tX��3E6�n�@	.��q����s+-��$O��R��9���i���h�L���҅�ԛX�z�m�n#_��ӽ��gM��CBÆ��V����3�|9V�,���N`x�JP,��jġK~�J�C�tA���>Hƕ:�OjK�+g�&��g_2�;�v1	6���9�r���5�E���d%�Q��6�8�*.K�?�U4���[���t����FH�F��}0�,���ѳVbK����[;T���A��J���A����L�u�k"�����t���:
C�j�}k�9jv���37.���W?�<�P���Y
���{X��A��G��?BҷXϳ�e<kO�K8�:H���¿��H�{/��������/�����s�]y�_��V�mvJ�o��I�7 ����p�ŧ��h�ӮHx0GK2i"��E��B�j���#�����y���
�j��s_�"�3��=�-�9��*Q��1F�T���B[�C������F�2�:I?�y��d��ԯy�Z�c^H���,V�1�n2� �+��&;i��l���9489���*����`�7�jܦ-�u�?���-�Ҏ?���d=�2%IN3���d���r��������.��K�if_h>�Ů��9���LG�__�]V���f&YU�����B��&rց��I d��cD�'j�{����{�Z�rlM����l��	V9��gR���:!�Vt��ˌ�u��o3��y ��m��v��v��dT}]�dkX�
�}	���#�׶TQ<�mQ����gt�(�h��AYUB�Y9�E����D-����r�IW@�����{Zebcm��-���|{���|}4�/�'�	�Ť�c��8�P%}�(�<����8[Z�Ϙ2�K�:#).�,ި���J)���id��K�Л����Tr+��$��O���O��䓏�^G�j�J9�]��0y���kl�P9��%U񇧏FeAe��J��QUY�et��o��G�Ys�, ��y��"�pz��o"�����8X=��T�\-tQt��wN�:��ϴu��S�`1y��+cj�G�0*�@Ý�.�!̼Z�fb�yhuh�qs��I�T���[�F+OL�<�vVH�x�ؖ�����;sfn� n�&s�����3LM���h�,^w� ���̸�{�Fnd ��>I�'�{�(��,2���0z(�Y/��a�o�路�[j@�*T	�v��uA1e_�k�s�<̅��x`=��u2�-�\�(X�1��o�"�x�S�Ȑ��N�T�<��x��E� t����������?Ãp��yY9�hI3@nx]1��{���haz��]~�\��J�}T��}_��QĚ�4�jE���.�z��b�?�Z���cH�-������f�Bs3c����D�����f H�� 0��u�\O�-���`ƽb������"�+�[�Q�:�9}����⚿-Pt�rU�v�E�amx���#*�_�^�K����U�l�o�չ ��+�O9n�X�q"�X��fo��������Yo��*��d�x�o�+$�-�[:@v���G�[�Vn_M?��L�;d�bb_#���h#?h�����	`
$TE�����i���B��{EC�-Jط�x(������E����&: Y�a i)�i��ʴ�f��~���-¼YE�5i�a}z���C�^U��J�)�i0(˝��ƫ��B�����F)��d1� ��x>�9���A�3z��"�����n�p�9�cE3��PL�M�P�*<�R"�_0ӟ��tm2�^�������>=��$���PDV�	���Rz��,ð���W����G�h\��Erȸ��<^Y��ݐ�ؗ1�;a�N���k����̨��Bt|�GyIS#0T)R�1�q�D�j���M81*����ĥj�������mƸ2 ^�S�.ZW�f�`o�=hi�MI�u�p��3_�6�lox��/�:���}Zb�s�l}B�Ɋ�ZO��hP�8�w�}����!�hq��T��/�@��`w���u��z.��w�mc'�b�<�v�VGeO���W�X�A�[��w�j5-ߢ1�ӕ��o`�t�F�Ƚ�F���+x���13Xz��+����VlNE�IR�>��-!�QM��� �����pr,V�.��<��n_�?{}��<N"N	r�Z�{���c�<�1���3��6��K����̆z� ��}5ٟ� �S�r"�E���,kaa��\z���O-�����~��Qk��;��@wj�^�1�6���N�� �G�R����K�u�;�fa���q@�,��Ǳ.:u*�n��3����<���h��q}��΋�O�U�|1���S���%�vXșYE�d�hVN��,��0�����z�f|���s�� J�홤rM?����à��0r*�S�'LH9�=g\
#��
0�0}�b,��k�� N��f�@���ǿ��j�a���HFiZĔ�n�|"�å�1ðt(��{0
U}�h0�5x�~�\U���"�	��\O���JP�	��,tUP;P���I̼JM�0`���r+
�����/���)�w��o?`5�b��K��z��4��D�_0D�lA��;����V@��?�!4�e���a��k��(S�W��8*]������w�l{��w7wȭu>�	C1�������������t�s&jˢ7�����6�	;F��;/�[e��Lr
���!ކ��ȩ|�~��@�X������3^56R/� ��*��Da��1@�%�s��W$u�h`\1 ?8�m��ڔ�Pf^���=d�
\�qX��xA=>�\	��nruʏJ
�V��y�c
��a�ǂ"kC��;﬇���=3�C��a+�Vc�ى��ġ��;�+E�Ì)>m��Nn�񣐺ۨ����r0Lt)��5���/�?���xd"��dl�Q	�R!o΋��r�ំ�+�Wgy�ş:�(#Zq�Å|��q��w�_��<�&c���w�"�ybpHiQ��+�Y�V�*A��
W�_y&��9�Iq�����`Fj�����H�Ů��8ni�8�S-k������r�����!j�w�qKWFf7�|?<�F)�  r���7���j3��1޷V+ ǖ�ˈ+4.;��m�+Z�w�>�]�}�_�^�@��z  ״9��0�.῎�ֹ�w�w�PP˒A�80{S�ϛ/�7o�ٳEY�r�
�%�^��݄Edc�v��#Ĉ[!�̵>W�>&<ؗ�t_�Ei�}�-��k��~3Č���~}o��e�;�:�0O�:H��������(]=�>~�p��+3��̙tj���pd=e�+j@{�RK)u���T�2������Hp9<<����c�p@���ʹ�l�%�<hPw�:-k�t�,I���i�����n5���
 �Y���GJtb���w��*�%�����M��D�c�Eq��l���b`@�d�6(brd�����B��nQD)�]Klv7�j�Lzl<�s-�D?$��[�����x)�s�=��$:�gf5&$��~��e�ly��~�!���[}BU�!q���A���$��>��T�d����-���,�^̭�Dw�vU��$�纻OxQ�/d$�ץ���w�X�@ɰ���n���AR�{D�9�lP �ћ���vN��ނ�7N�F�w�&$�e�
���K�$f��֤�l7&�������&�yƾv)��z�����#*�Fc��@ /H�#�D�Z��k��X����^�g��q2]2�����Y�Y��?��p�̌��]Z��)�����eL�F����
?2�_HZ���Z*)��J��Y8��i**i-�U���.��1�a���Hߤ�^�z_f���~��O$��P��z1wQ��qw�`�z �3gXc��/'#��^L�A�gR��_ݧ	�(�+�:'�5/偶N*0�p��W��<dM�C����i&ι�g0��ѩ�x��!���"b�۲a����U��5�rNɝ�/��E��u���N�Z_��Cg��d{(�ݐ{k�mձ����ϝ��bP�*��e��B6>]���F��l�� ��֚�ȑ��`o�I�V���K`7Д��jj�T	�Wg�?_C�W���͜.�!A�8�dg��[�����^��2���	��Tߝ�}�8�#�{�9�y��n5͜���K�W�u����{�0�@����ڋ�e��Y�p&�,o�;,Q?٫���}p@�A���y�*!=
̡Y��.:�x*��1kN�^K��ާ�Ar�o�v�����KJ�ܷV	0C���,�8��B�hô�N��z�Ox�Q@�,���~�8ؓy�aN
�ٟ�=����xi��B�������!��t	x�g���U�ߌþ^�n��q��ϱ��k��ٙI;W���j���Tz['�/n���K�+��[�Bc���R/�vZ�T��1X9�݉�9i�nm����pL����������5W�v��|�������]4f�Hl��a�?|�tx�� 	^��z�	���b���y���,����~�N�5)�ţ��̮�>��><�~v��+]�i~ �j8�aGHzkٕR�Y�'�bN��>b���%��ޕ.l��i`dýr�%1w��Up�`��~�C��ߛU���MT4�1T�y����$��n�������9�i"����a#͛p��d�����=p�Y�%:�J�	���6��Q��g�*�I�����9]�������kA�%^�Vݨ�*<N�j�J��Hi�5��s�4�
�b��ˠ�$k�?�X�e�J��$҉�E`�2�y镋�M�)E������oMk�h�d{3hH F�U9��>_�ʟ�a�a�lV�m3�����o��|5AQ�"���Y��4�rm�}OW����R�� �}��Y�?��֍sԩ����:��Il�*�x?�j��n��Ї1-2����DώK��A�#�n�I�[_uJ�6e�m�3�lA�tcTYxV��~�p�Nkm6�<�����霶IH61]�ʆ��w���{�>�ʆ�%V�B)��5�>�?�g���P�O�]��EO/P����˧D:�Ook�����۾�sT�l\7�6lb ��[?��̃�}�z
�F\�<�������� ��5�CN8D�,�t��E&)G��EY��3�"1�%��֣�?����~N��9!��z� ��%lMM}]ƛ>Z��Թ�A]���?�[�e��#:�IW�����`�s[�%ܩ0:�Dx��Bk@,���k�(�^z##_��nox=��T��S�
��	��ǂU����ʇ��'K�s ��
�F��s�Es�<��$0���DN��騷E�'�ȁ��Cz�\0!���7?�;�K��q�A{xcw��u=���	��>�cM�1J���	_N%v����l�`����coԑ�0��c �h�%W�R�	��VP/��96Z����w X�YD��;�#!L�0Wy��	�1[W�^,h�����$q�Bj�Y��$��ҢP�!�W�)���+_�H01"�������8�,����Š�H���D.8G|���+�&a{@U��mQ��G�}�%�+I�Q���l��e�\9$Q����p=03�U|􁌁T�;��=�Q&��Qi�g�Inm�e^5FȍKt�������w�};�������ß
�_�b���[�)�@��͍�Jք�N��A�j�z�:DֆT��W7�V\��&���v�����>����^w�X�sV�=N��J�'�em�p�
�ʍ󖂛
�٤�aq.�(��@'�w<��զ��Si?��| %ˀft�.۱��"��G����7�P\@�k��
K~���cѩ�b����I&�\��.UiK�-t�Ԍ��͑0���x%�#�e՚�����Z)�Z�(]�j���y�|ˀĻJG6W%�{� 8Û���l$���&W�MB	�~7����c���-̕\?�h����O�2���Wo�~�2�*K{�m?6t���t� ZVb1�>I��c�^+W��H7$���'V�b.�� oa��+c�U}�Y��]�b���f]�^ ��/��l�sҡ$�`�x��	s����F
[ߖ��z�\���-I��*�w��w�V�c:����䶡�+�A��1B�U������M��+�& n��٣s3�s��E�I���B�2�5̾%9���ҹD�^H����UI`+�}ι�O�QGx�Dq��{"��U�B��u�5ƚ��d�?Y��K5d^lS:B��0���2�; 2F���� �F��ʱc b�����5O�]�qe�b �.(�W��.c�b����<�}�V	�nDe�(Q˚���m9�Cϡ � �]��
��z��,�H����Gz��&D���)E�گ����QX�^ $Z���S�Sbb�bL�}���cM|#�W�����&h��+Q�!//|�k=ߠ������%�F�!�8�}�XL�?z�+8�,����@Ms꿎ߚ�,&��Lc>qB �]ta =m��6ɐ����y��?��8�_����٦��[hȰ����k
�d0O;;��v�ϗ_�Ftx��%���3��d�:�5D��Z1[p��Xj��0�Y��1�^��R��d�k�ScAGkOu/EN|4�xU���e���~�A@�+���n�i/��6����D]�[^�́��ef�oy>�Y�7��̌�1
�.�&XOM�#���-��38�2�����䙉�� ��I�U$��d �pBĚ���
:�&�|�Y ���+J�^�g"�+�J�l ��%�)ݲ:���m�5�kޤeb�0e%ę�-���{���5���5���(`�
]����.�$��>�ےϠ>o�����?�4ź+��U�X���2$�4�������{'�l��s���.H�}Vmd3Ϩ�>��R֩ ����p�Z*��lF?����eh�%/��&7^�/YD�&��'���u�����jv�<��5��=���?�^�Y�P������︎T�����MZ�m�b/�����=�%D�q���)�<��m�ǱY������3�ܐ�û���l[�&�����M�~
���Dެ�����2��/��W�)��R;��`���� ��9����$.����^c9F��D�q�K_�&��a��A�wLwݤ�Sý�LO/o!? &�W6�
?�v.f҂iuVQm[��-���5Q�8��*.�į�I�
b՚�%�7~JSqE�Y�_��'����B�Z��mu#�$�xt�?�a�W��Xv���*��P�Z5�7"�˛��;
�X�	�k�_7����v�¢��/�aJ%�h�
��f1@����ו��x�����xĵ�9~�.����F��*�Z�Y�8���[BtWguw�b��S���QTo����a՟���}�$�����ZJ��H�78�)(oX��
�}����<�*�صH�sp4KE����Ϊ����qw��]����L�-;�����^m3��+_z�@���QR��ǩ�Z4�٫��j��ɩ���Cq�Z�H1�9����sKm%�XB��9�=��\��ݶ�]�(�l�
c��a-R[qy�$����&��7�=~�z�-N��L?�:�xq{��B!A'�+�)�Vӽ[\����b��i1eV�&Ȕ��a(�_j�l��+�t�F��g��6V�vX���C�r�7�a�Ũ��l����L�K�t�P���Fˁ�&��3I%s$ h���qY��\|l���s�Ny���5Aܗ-)\�Bީ��86�/d�o��������r0�{���۱'�4T-�}��g�??E1O2��(6#Zw�C�a����EHuT|�%��_�Ǜg��
cu�Go��4/���/^FKv*)�$�����)�rWk3plqH�����ԻR?s�~����+���D�|�?���bb�y�u�ӆ�D����
Jaʳ���j�o{�^�U�H����5/H&�+���|�hI�	�R�C��X���
�a�wx�`t ������w#�<�l��z�Ҏ7x\���ڹ/B|��&�f�c66�W�Y�dq����;O�tDO�
fP3�a��K�Q� ��y����:@2�U�/홅����LsU�ؐ�C�]n�-=���I
�D�_�J8�Ɗ���|��w���1qi��A��]�1��77�#�/�*W��6+>^]yқ���r

��X�]9�&��� ʹ���0E$��Tї�p"���C��Ǫ�:/��$�nڬ�U����V�ײ�Y�271�}8p$3?un��72�1�	x�Τ��f�v������_%@(6U�
�wm���v��ߜʟ�=�������uo��wZ� �����L��ħ��H��"�:j��`E�����g���͠r�:r�Y��o����a*��5�t�OQl�aa������HI�7�9u4�ޫ!��
Nɗ.�4��f����1 �bxF�f�eK��Ľ���4�(�	�K�"Q�çA�S�r���@��-D5�t�s��� ��`^�nY0��PK:;˂Y����B��_!�5u���Ɯ�^14���+>�[�1����1�Q��u����%y�z.��Jnp͑f�&6	�n��Ν���W�;�L����Ʒ�}|���W�bK����W*�$�l��3j"U��)\e���Ɨ�l��h$�N�����M�K,��촏��\na_=I�������8�c��y%���acL�m�y�^����iD�&�x3��?!��wiW�<0�Di��&��,ew�Q�#[���"�	BQb �R�~�p8U6�Gǳ-����������H�	-lY%��#�z;z􏍑�+��D����c����\�A�=	3��+�!�j:@��+�pr@��b�8%+��	$�u�(��G�y$QZ>�H@u�6 ����T���̣5�U/AR�3�ƺ�m��տ׼Ux|�o���//�7��BE��e	�@f{�[($++�`�R,@�Um�F�E�j�i(Y���f����̓��tqQx�����n�)�a�,�Ɉk��N�n��ex1����I>d�:�	����	l����ٞ>���`�g�+�~N)<���z�q�տ,�Nĉ�C��0�2�=/Z�r��R��0�@+	v�[�%���*����ݦ(K��ͯ����������MC��H�N)�<�T��!DB�|?�j��7��@���נ�'��l���ga��h�#ܛ�N֢�ZW�J�FR1&�b��#%"~#ٸ�gK~�0��GTAC�Wl۴��	}�P����00�����0U�P�����mī$! ��i�i��WS��PX�>VG�l�X#@a���{�L3J��>��w�0G�4�f���zx��_a��h�R1��<��#Z�j+����Pz�Gr�}�6s�����8���q�$d������0��*
����1����.�Kdp-J���A(�ȉj��G4�}�ſ �Fݧ0��6	Jj�������	[�q+�lYN��%~�	j�v�>]��z���f�@%s)������&��s��Y�(7^��O�3�U�tA}P�QO0?�``�����?�)#H(&�1���lz�C\V/]t�����!�J��
�A��wS{���:���
�8��*$�z�]����K��x�����!����7���b[����]��\�_!^Z[ ����{j���d�+�`���b��O��q�I�)s��_���"�C�6��2�y��#��*&��u��(53r���U� �\V�a�/~���[����!�����x]�-e�o=&��ό۟t����%����g�M^Wb[̑Aoh���xc����N�4��i��9ʐH*�%�'�5ٱI9�0��U=�����)��7���[��abY��0��ֹ<r��!��]V+�Z���2_>��&�k&9��u���x�W&U��U���e��"\�;�ݫ��ĸ�U�򍊪�;py��f�_� ��?���<ߐ�
���E䇲iI�Y�/X�\"�[j�h]ϱX$1hM���
]P/M����M���ZSg-�QQ��7�nq���B��#G�L���.�n
�eqB��3`�:�5�& �yϜL��p:��t�j��pm�-4�x w�5a��+ȭE�5l�@	�q��np?�Np������Ky���"�=�5�U�d;�f��9�P�ʀ���:fK[0���
���?��+-�:�����o��vٛstt`��&���L1�}��1R��`���7q�A�ͷ��geXԓ:3���9���tS2/��6�h�N�|�2렏����6HuI���uJ��~�<�?�nWqA����ф��nm�$�������Σ
��G_�>x�)����+.:"��yi�K ��G	���w�J�׸ ��p�p>�X�c�(r����b�
1u8 ��8U�?�GF��lN�R�'�D��hܱ�>]���~ݖ���1����Y�� �d��h��I�Z0/ٌ�����*/� �a�)�L��Mg�y�9����㳯��p�kc�$�����z@�����$}ިX��� ����T{pp.c�%�O�4�9�8���6g���8bF��]����Ǒ�L9c����a���-�������4��;O�8�V_�r��ր�n�^Q�|�)՘�C���c��5�z�+k������G��Ł�hժ�\j?����M�vuԶ�p��"��C�¼8�;���c	�ml`�N� E�!�9�na-.��Y$(�hח���[�蒱GVeI��ƊϷq�TNk�z:_�/ԣ{PZ�"C�h`-t���P�''c��$���{V\�`5�}�]����;��2�b��ѤB8���&K�ܽ<e���Ϥ�C�J�;F����ED�Y9m9���ƍf��8f��t�9�Q��uW�ا�}A(�ь�,���f��� ��(KR��w���	���/�5B�
{-�XƠI�-X3��S�&�E�9�/��OV��Yj-����<|����K"y�ٜ��J2�8���OC�(���A���/�@�a�_��r��.F���W�A�/�@�2���"�a�m����h�� �N���\�̉��CN0��PA�K��(�*=���&Vi��p�����LM5&W5�%��ub�������><�i�;@�*�L�,�%h��S�44��℀���K� �MT�w����v�_�[��oʱ��+�|��忚wQo��tk�����W,9w)ƽ/�j��ϔWD/򇁧�E{�*���]��Qv@�i�{��N����a�IO��BAS���%V�T��ڠfyOq��\#ݐa�!k�TJeb�<�� r�^�&($^�vo�G��.�T�r\�ш���s|�����!՘ٰf��Yv�̝�'�|�Uc�}�V���z���J��#
j?6��fﲘ�Ge'~�NoY5F�㣃�Li��oj�����(BD+�\Sc5����qT�s�CZ�vlrv�La	ˏs�{%���H�7L&R�?�X_Zp��uҞ͜��CM�s�.�^%��[�6dgʈdן�Ԥ�]�0�_��Mu�
t��N�B��zjo�D>��y��`^�Yokݴ��͞��6��k[�y)�oR�~iƥ�6Z��$#�r�� ��x�DU<��
�H��]9�S�.r]mTL���3���;c��;`��~�>�]���JBGF/�'��h��piS~�4 f�(VK��"`�|����0��2�wP:��)��y��v*�~�u12i��(��.M�>����k�E,.�.һ�g,{V�!�&��e5���������?X��7�\��=rRT9���NӺv��U��,�r.�NBedX�C;/r�CS&6�]�	�>�Q$Cp�D�|��eL�ez��L2��0�j'��-���c�'VN�a����/oOy9�	5yu0�=l6��/[J�j��N'��GS�����MZ��<(��H�g!�IU��Vo�mo-���Gd�?Έbv���fXOT��j�I�9;��!~���ݑò��F��q�D�Q���+WyGmm ��-n�+#�j/0����f����_ ��@W�봻�<�9���  z���P�5�:�!;�eۭ�	T��I8�0��2�U�5]���.E��j� ��<�(�le���Ӫ�{�RK�(	��J� �˟��[Y?���6����P��RQ/0����@N�2��pLf��
;���q4��RR0�/f��O��6p�����70�ۮ�y�SP��4�-Yp����l:_jɅh�J��%(RYy�y����# �����hιE����ݷ0G	ʂ�D��L,j�-bw�^vB��ȞZ�l��m���g��}�Z��{yx�L7����:�\��P�ɲF5�X����׶$��E�O��kh+� �9����>�,���p�Bl��f���>�pG�B�����Cׂ��i��`u�c��1��L��h�$躽�}u$�aKk�3�K��)�ӎ�Y��K8���ß��z�NTU�DO:}B?yی�	���ȋ�*B��#���t+r���k������y>"c3�&?�Y�r�1�7NmF|	63���S�i��`�W�:t���Zlj�3��t��u�h���IL�xە�s�c��Φ]UT:�u�ʶT �����_���̩���0�A�Eo��d�Ӭ�� ���W(>���|�hE�0q,5�;�t�QKD��\�@��M��N�=��� ����'��2��]����a�#��~@ I�a`��ŗR�V��5՞�J����qb�N%�(N?c�	����K���W>B]"���i#�W�?�ߧ��R��n#��WCC��-�������^����\��;�cp8�D[�ψ�s�a�b7�m�G�)(�8e���"ܝ~I!i�E�mnZM0z�0RG�Q;���74�N�}�Y��Ӯ�}�1�24T?��ڤm#�Ϡ�ZXs�q��=ߐ?8��� }ɥ���������7�QV��ύ���9R�H[죆b-d����ʹ������1`q������[��y{�������*,_�*�!V����)j���`�s�J�y�FO@S�Mdl�D1���� ��-Әc���:\�j\��3͒b��Z�L�Ͳ�/���\G�����V������:TB꣧�m�s�d���p�����sp�N�cJ��#��MJ�ޛ[�~2ws�ъƠd������hz<��e�U�2��J��L<:�cEs�����o�k�QSE��R˯.��Kx�P�v"��,r���ȥJ�ˬ����ǵo�-�\D��g۶ I�{�Y ��%� -W�$�g}�a�\JS��:���N�p2]�+Y�X2	��v&���"1�������
�R�����u��\ٜ[}qKG����V����5��7��z��:�)��}��.9�0"�?����2p�g~�<ߚ��-9v7�c����P��fQt-�t���Ak���1O~rI�Jpdr���J����.�2�阢�d;:2�@����WY��$��|j�uB���>�o�@������=��r�l"-U�k�!���MPS��NPs�
�2�1aWٔ<B:{�h�*�\�?p�{*��&~��Jפ��{�u��\R�p��Oh�����ǚ�Mi�#��Е�%���P}t�iY�̎l�$!����$�GJOs	�#?�7*Rc�[��χu���pT�?q��g5�V��2�J��/������Ą9�F ��a����jm�Q(�)���{p;<�޶��YƼ<����v����3�L�`gK���#	7�C���
/A��{#���
IA"�R�$�h$c	DЂ�Y� ��\� Z����9��p�hR���aZe��,�f2~(�B@g95-�����'����gl� \T8�b;�xk��Jik�Z�F}�;�ѵ3�� 9�c�TbV!G�[ �=##6�SUPГL����!N&H���M�S���uq��	7
�~��K%&Z	n'�؎]D�R����05�^�{�^�i��W�w2.�u��0��3��&������&L�����1Rcu�K���Q�90�<c����U����y}q�Q`���s�8t1���Jq�<c��F���_K1W���G�i)D�>�:�G( h3���j��LDC"{�9P��
���J:T��6wޘ>�WɗF��E�N����l"Y�~��+�d8���8W
(d�KP�ۚ��8�&�Un���sfР��hB��8������*����ٚ�&�gN��`���v�M�
����x���B%Iwy=��ך
;����f�z�0��F~�]Zy��Sf�kz�H���75���;��S����m�-kH��~�]�e��B}SFy{X�Eٻ�V](fְG�8O��\����M�����.�`�7HꨡE=�'S]�^���ݜ�h�is<��gbi�v,ܣ��������M� �j2�-�I�Ǘ�B?�*��j�y=�8Ě�7wYg�;������A�nF���G�7`��k����������3�Y���:�_��`\n �_m����ņ�&�����9J����� ��A��#��k)+.�<9寇��&��sP��v�ܻ���O��J����\��ۏ>���ǰ.p��C-5m�\TicFlU*�*���a����V���'�зq�&�2g���!�dZ[���|	��g�2:yVq�
,��E^�S0=�x�Rb#J��D�~&�-Q�T숯��B��.���{En����	���4�we��z^]|���?�c��>�ӎ��տ��3ƂU�j;	Fb/�}/�ݏ��ci�*�)6��)S2���k�Q�ސ� �U$�[}}ҙ$��-�>�3�ʧ��须�ܧ&��/<��4�7���{~��E�P����ۀ�b*�E��d�M�fJ3���ّN�9�@�75�o�6	�1m�-✫r��Z�[p��=y�U���]�aXw�К��H�b�7��?y�=Q95h���`[��&�@V� ,���m��n0�ȹ��coz� �IS���z�2�D�"�������w�����ӣ�ǌ)=V�?��nx�Zn,���ȐU���ue�CTwXY���R�>��kp&����Z�Y�ŕ����'�+ł\�ސ󃔴WW�%Y�Ⱥ����	X�W��w�xz����`A���?�懇�1fG.d�2K���So���F4í/J�>Ӵ�S��W�yn���&�����>��Y�YI�J�|�d�b:�hj�l �9�oNh�<j��!��`gew�1�����/Q|�"ٞ��镛��n��S���@y
,�,9�����������Jt�֐��t�o6�[���4YN�  D�b��u�������m��
�U�x;ˠ|��h�I�J�7<Q�O	���'r�J�!��IE�[��� ��Kn�"��3�J�o�a��Et�(Q�B��3�6p���O`%��dI�m~�����$C$G2s3�����c���O�S�p�ú�>i|����n����8W/9�:1���(��2����s�T���S��)����N�ǵ�m']�x�/Vc��][��i�b��m���,���|��ClN�O�bu3V��]�a1l�IҒ:�5"���n�)���Ϩ"��j���1>HC7���k�E熃�ޖ���H���sc�u�R:R��^_�v��㶀��m�X��YE��Ց�X�b��F��^���@�/ޡ
U:G_/�p���S���i��v�.�i�FM�I��:��@���5�9�cl��2N	�*g_��і�M>[,�瘅��S��'�q:����wO`�5b�o�y��`�䜖�e��K�%nr /k�Z�g;��E��l���R��zgy���l�g�՞��ޣ��:HRm0����Y��]:�������%�xuPX��'r[�7f�����H��S���g��ho���3)v����k.��q�.�B�{�_��JQ1{7���ud˨V�̳p� 앮]�̔��V)�����/A�NS�
��B�T��OJ?�ա�j-#lN�H���P�:;���g���s�I�[�����-?�2""odGnTy�� ?��F�����?�}U�xza��c߆�u\�Kc�u�`�RR�ָ�U?�����%t��+���h��>�7�����U�ɺ����|�1p�Pgo�Y�%d-�~˯:G��dM��mfqh^�����&~�,�V�T�/�w��ҪZ�)�N�B�������\0�#9��T }C��l�I��'��+��4ک����d�l�=Q��TV���X(	��6���,��Q���3�`��Ԉu�WY��@�̜i�&C^al�G@a���`�Eu����y�'����;~�f���y�8�1A�;���Th5���b����1>R��n��en�ǾШa.�+t��:s���Z�����/�@|i�b���+��UY��-o��a��ӣ&�H�eN5���׿g�2ޫ�P�ލ�dʤQ�_������0�����E�$S�Y?C�-�ɲ�ɹ���?G�
l�:����V��D6������u�'8�7�`��[_�Kzsٸ<v�xS{��a�*3bi[,�:�;`�|�`��L� ���m�_�G�1<�=�-�;3��
�X�l��������^�j�G�I�Y���K��_�Ok	�)�q���x�(����/�i*�\���y�i��_3���C��y8.�|p�B6���R�������+�����>r��Q��C�K$dc�&H���\�h��o�C^a�9K�;*�6��($���W�I�aH�팂\��D>	�Ѝ�j�b\����(�NZ�`�3��i�	&
ۛ�iب��d.G�#��4����;|7��D�bGhP4�m਻�irt_���Iߠ����P*1�BMӕ��>.`��:X��D��l�
��S7���焩�u��#�wɉRw�/�$XɈ<��V�U�?����C�f@l;��>�9|��Pb��+m����h`[5?u���+��1n��>w����ٓVJ�k��c�T���ֈ�| 䵎jJ� ��3�ᇯ�x=�bޠm�GW�Ԋ�Rͧk�V�eƈIG\������ߎ�[�^�!��dXm�7�E6[��u����	N�[���J=�'���s�9ԳƳ8���)�5<f��P�4W��mlE\K �2N��W��m2F��T����dk,���܎S��(�*td�5���*��q `��?ABЦ�}�����[V#���6L8a�[T%�ȕo��!Z Љ�X:<�R6��T� z�Ø�O$�z=�>����@o�� �(�aa�H���X��HL�Ƞ�X����.��vB����l������_oό�X�O��Q�< 7"�fmi���e/���H�!����7���Y�������.� >��Zv�Le:K���r��14��TY�4Ww��\|�i��94X�~�k���k����{�Y������������w���_ۯ`�+�%7�5��0)5�f�b�<zB��%����<H�cZ+��	�fsd��W��g��X���;��H�r�9�9D�����jo(�,2�o��(e�Þ���@�*d�z&��/~���/��o�a��c�6X�������d�r�Gk�:�i��,$8����F󔰨פOc�NX%c�qu2��J�:�A���?�|<�����ߏ݋�8/�N]�Lԋ���/�1?�
�`��{�a�N�_,�
)��ND���5����pg��H�|�~�@�-7Y�xG�H�����*���8�$�F�z�`�c�Rc��Y�$ضD�c�E%1�/A��Sl�!��Ӳ���݂�9�rXn(��W�b��n�E$�b7nQ��:��s?ς�nG J.�nc����ig��
]�Z��b�z1�H�dx�>agO�x��}z������uSY�?��A��a�ct�#>�aTuw��%(�	��q нJą��'�}�����\�ܗ�pZ\ym6;?̲��Ec����=^�-.�L%�J1-Qz�����c�QZ����V��Ϭ�<N�(5����Ӏ�:#�|�#�nq�����)�س�c����dc�S`��.9��U�S���X d߱�SEo\B��	�:��LU_틧�n̡��
k��a�d��X�ӓ��@��˧B�$-y���E-�8����ś�ߤ��Qr�AҨVG�ʽ��6�1��^���z���p6Α1�#�|ϣ��з���>�I<��vޏ/ X�|�$����7"���0`��Ou�{��{���5w8��"vK�<�;��a�L�?2��z��2G/��������2d�a��=`!~��Y0�<�DGz��᝟F';2ұM����{I�Xq�ƥ:֙t�M|�<N�[� ��%�4~�qDH����� -�]�<�45%����H����;τ�g4 �Yؔ]�k��*z��u��ǹ�5�N@a��[IaB�3)g
�zD\y���ۑMQ]�d&W��<����2c�
�6<��wC,��]�w���"K˅���J��N�~:?lhQP��'������~��g��F�����j��eǔ<�#�A�:��ә*��V��p�)�J[x6^k��zny���81��*�x��2�wbu��)��$�*8���̡]�5x�Sc�~���nW�k'F Q'��ޚ����Cjk ,�]�xX���Q�c�FфJ3��m�J��@Q��)Y���|�$\�Je�"��w��Q)�wK�dS"d�!��O�n�;0�k�e0W��>^4�ܾ�b���mev�R`���f�A�׫�řG�o�����0�qU�7�D�a�k�nk5��ɑ�rܱ1�1�#to��j���vو]JoZh�#�|#.�ؗp�\���X�H"ɷ�xx|�_�gL�����p��_��I`�"?��ǥP�qLv��mT��8Q�D2�}o6qWr�֐ՅF�h��8�5A�
	�L&w�	{FIn��Eֈ}�p@7]yBq�!N;�q���1l�z�3,^�X�oj�N86&�gX��G���D"U��*!;,�_��S�m�6�ẓ�A��wgr�����*������i*j�V��:�k&+c��!'�=�: o��rc��j��F"3Y��h������=�	��lC�f�u��A������7�����4��}�H�q�)�El���5�n�w��w�n��4K,,�|��3F��(�g���OJd ͋���p�w�&���'�?%oض��m�1�>~I��4���i�h�Y�57y��?�5~�T̩6������E�����F����7_�`���X\��/���@S ���/��-�5N�8��s����!g�_�Z��[@��i�3���؀��Z�^ ��_!<!τ�"˶u	��V 0!�f/�_���}`�ѦG�:��7�K'�m`��ݝ&w��%��{� �	��}���3���{��,J�t��؟ˀ�悥M�j'�+�(��� �$I�y��?��T�S�M�;`�d_�ZJ+޶�!�``�?�۱|��t�1ǭ%��T?�'5������,�j������A盨�
�:�������Vsj�~d0��jr�6��������'ݠu��<gM�;�4�: 0�ҕ�хER���vK���w�X��!���mzs�(Ov$Զ�D `�81g����ف����y|IuW���ه*j�|c;�7h�gPW����.t�WZ��]���W
<�b8*� ؖƬ,11�S�t1���X́��8�f /�(�XR�SgFta��bp+�K��S(��$&���(s���'N�nwC}S@[A~뺠��)��g��wX�
��ӑ�	�rt=\��ys�����Sa=�qQ����EI:GqSk�S��I���^@vy�ˌY�*�`���o�3?�� �ͮ���;�΍.�2��F��_k	nz⬒�W4��FQ?x��	h���t� ��[Щ2`F���ٚ`rv�gT�Zpe�b�GzO��?��ߒ�D���-��V��4��`���CΌ�IcvV&� ͗��]Yw�a����	��C��v�(��2�yXM^�ad��Z��4��.�}��zX����_D!�#�F]��qj8�_54D����p�@"{�ʓ�Փ$u M�P�����@��y �]��۵��I�᪱>��v�\	v2uW�Z���bl�ET(�9�ց���G�h�m���tň+�f��o�Ѿ!�5����i�ϒ��a��#��/+��8�_2�bU&X��w/Υ�딥�Z�O˛���9f'-�5�8����T�P_��!�*dK�{�V	P6�2D�1��x�mg}���y�`8:�W�Й.G��JT�q?,]6�/�jQ9�6O0��T:��1E�w���v7E�	��_����[TdM62)�p�����O2d��s��Č����I�I�N��Fc��D����F]b�6�Ɛ�ǚ6�Ħ��P�:�����U��@�pd"J��(ǅ��f�=3`��t2�
(G\��:�+���ɲY ^�#���8��/pi��lh��Ma�Q��\�5Μ��s\
�;O�5����4���{����B�v}B�f<M���Xחڂ���G��Kf��QI8e�_F !V#��/�>�D���}������Şm�bnşʪ����o'�n�R,�In�$H����HKFL�Q�@�����N�/1z�3T �K���j�ܮxK��!~�g+h[Ļ��ʷF,�:�ݰjy��󘰐�9/s�B��)WR�����kÎ��@������u��?���I�q��`����h&�K�����.�iO+��`
'6*߀&@*�Mwъ���Z�g�])~lt�$�}����Б\�B����m����0���b<ᰳ �):q|�� �c5� �J�}�� !ల#h|���6�D:C�VEi׃���pW+��#��*>�M�=4��<�e�V%?_d�ڕq�T��������/ƭ[';:�G���SgG|����轸�7>ˏ:9�j� UD2j�M@u��}�7���$ɖZ�f����p��(/Rn�ٗ�PF"��}h_�3��|6&�}��౮����4~��>&yNu�}�s�lA��
��Wk`f�8���n����`�&5'��.���,�N�
+�?}p��c1��\9zv&����I�S/�95lxa2���m:�5�:���aYu��Ow��cX6�@;�$�k�V:k�r2�ӐD��5U�o���P���}ǋ������� ��	�f�n����`���6�tۥ��n�Ovu<sW��(�sqR�jK�(}�Hz��^+��[F��V���YIdj9��A�K2ɝ<*�>UNq��I�A���;V(�c���t���]�[��mໃ�@�E1_c"��r]5�0�]|�0כ�j	ch�&��/��5t~���'B�d03�2��]M��Bo�w���W�Y��򳿟]�'��k���[�ӜN7Ѥx�Z��p�ש�Ƈ�����^Yl�C��.�� ���F�5l@�f��y�ަ�8~���.mwSh�Ir,�Cɛ��t��#��T����y(<����z����?$�B���<A<]��V�#��t���J���Z����,�\$����Ur��1���W}Yj$o"P�7|z�$�F� r�W\6���� ��lC��W��]��<!�e�H😷biõ��4{iE��Y�}�X�vp}^ۜ�6q2�t�? G�����*O��*^�3.���d}���$������>���M(��C�Q�`0!�g�0�.�ר�CEբ �Eo�o�҂�3����MP���쿎Q?IZ���vh-l&M9�O�@ƚ�F���M7jU�a_E�D��/��V}A��^t=���L���?�(/e��F%@͍�� M����-��p}'�)f����ɢN^QKT;RKVPk����8ײ�>xol^7 Z�P�	冘2��v���[1��	ϲ�B�n�6��E:�m�g�ݡj�:a_O~�LI��	�ǋ�� "?IAm�Ę?3
�6�� pi,�wZ��L<�������Ջ�b��0�P�
��2ƭ�)���$���i[���1��*�2�8JM�a&i��d��V����-t��s>{4�2Ez������n���J�O��.��
�7�*
i�F�qЏ@�S��霥5;���-cF���o@��l=YJd%��G��!��4�Z�[_9{��5�W���"��@;�m��r >%�XH�����\Xi�]�6�(��s�x0V�M�zԇ�@b̧�h��>�DU�rIq5Py�3dM�����2�o��!_�l�cN���j��Z� �NI=�l��>�{�HNu��a=��!"{�ׂ�9,�4�ХZ�VN����ȼx~.$R^���U(��v�g����ʼ�d�<��6���g ��YEf�ԏ�;�B1���69K_}��D1�=�TK�K����if�ϫur�U�8bt`t=8J�hR����T;X'�=��C�|��F�<-�0��z��ӛ��=�IV��{�H���$�����g�冨�|�"�cH����{����h��Sj�к�5�J�͊�qpg�TE��>��C(4G�Z�C�dr�8��ȴ6�1�ī1�\�3v�j&��=ܤd��8TM�r�ֻ��PR��;{#���L|F���G�1��T:19��9W�Ƣ�z!�c�+�P9Dĭ$7tf�K��td�����D�RS��`�^�?��$\WKzɻ���*�����s 䊵����	�UE�m�M{+m{�����"qxF����@ �m���**j�FJ�H��2u����WV�/���@:ʪ�%���dR ���mC��Bq'`y�1�e]�ܫ�_�A$����4<����,vj���iP<O�U崌)��N�����s��J>6����;�®��X}��[J���RҚ^�x�_�TM+����l^v�$�C�c
��!�[b�+�d�]a����P�O�(�z:�C��9Al;�|�'�7�%�V�
���ط(r�{��p�	yY'j\+�V�����Ѐ���yM��t۳����;�-�Rt�BS��;���#Nunrm�;΄�4m(id�s�6hE��_� ���9g\�z��������D]�Q�T��ü��1��-3y'2�xmBE�k��NF�S��>o<*�3�p��c�)A��N�dh���{��;���
��߱U�}�0+6������.k��m)w8�.���|
�d���k�����\��w�!�f^�Fnt�[�ƛ��0UW*���aX�@tx� Ŗ�ƮH�@�s�N�����>[>���\��(pR�� ���;���A �"�����D�&z᭮ 5�]&3R��ԩ�4�^)� {)s�.:��/�g ��_��1g���Z��X�>J
�ɳ���x�|���`��~�0]aj����)�\���[*:-W��2R9B��Rft�ds�i6ʃ1�'��WK��b�#�J!&���g���ؑ]W�c>�_g"��Gl��=��ح]4�r~.Q�������έ���x��nkr�8ֹ#�D�U�HH�ѹ>DQw(���5]2R�h�-"D����D��$!Y7�kAq��m-�O��a-`�#���m�,@­� s<�|!�
>J1W/�(�h�=�����}ay�p����Rďϼse��H/g�\�/j�e/���&�ԁn�(�m.{vX~=�0��BTy����N��x68���s�2��ckO��;�h��]���AyAmw�����#��'X�S�9�lsU�Pι��C��3����$��ؐ��0v�������W����oϻ���L��_[�[���)�-��?�ě0?���3�	hǽ��N`���x��H���3�:=���i�������uX�Xj�k�Fqc��P�z(�*�=�����eiG��8:J�(�"��j��-��lu��H�BFU��a��,��h�;{Z\���`�(�$�ͣ�hp����~Sb�'-�ti��dU# h@�YU^nZ~�0ng�
�e��������2S���s�"�[��-�mtV|��&[�j�r�Q�OF�R/�eW~7e��~|:���n�^�/��͐4�5X�6ك<�����*�`�j5Q1{�F�گ�����uۅm^�tW~����Uj'�k�D��ҹ�-�^��B��s擁Wq'���3>`���͸��eySū�<�W�7�~b����'����X�����E���c�~�{D<���<����	�b���F���4wQd�Df���-��R�{s���6��Ct$)�3~�M�+M��ᘟ�B�#�N���J��x�.Ga.!�-�� >�P�*s
c:�=�z��e�B��v��I�e-^��|�~	����K��u��sP��� �C����fz{9D� y�jq��腋��c?���Z���U�᫤��X6���>A��U��)���R�l�[Zzx�C���yBZq��~^<GoQo#�������#Su�ߍm{���9�_X��1��?,������y6y0P�'|(PҪ�~��J���cڌ>����(�����|�[P�}���l��V3K�>T��{8�9�#�zKMɥ��ؕ'6�Y;��w����	2QAL+�p�?M3%���HC"]	Ѷ��e=�p�PH��2	1N����}��~"��"X>��k%9�v��N�ܶ�Dzs��ȋ��n�A)R�������{J䊈�CQ�s�������.5��]���*���Ρf�b��*��Z��`ѓ.Tc�H e&;"��-�T���j�`����2r@���o�g�L���d�>8��KD�ȐN�(s$_'^�O�6{�8�*�ą~h7�9㥪������S�C��&��v�Fq39�;#k�F2�4̠��5ՆV��D�NwZ�,#�Yg�v�zs��CW(�J��"��99C������s��?@jIn�5n��G�b���&(΁�{M�(˕W��|Q���kw���6��7U�y���\\��e�8�����7#G��T��_�b��v��	�S,O��
�&�-W���e$lU��2A�`�2xe�S|�o�}F��ې��>�ǡx��?��As&�ꫣ��dK����Ƣ{>���D l4q��VhC��CKz����?*��5Ҭ)�I���b�������[7��ފk�n���nD˩�&x�\��޵��캾q�%9�*�j�!}�r�<{���{�M���Ҧ��a�.P���-S�xA�w�%Dg�/�T�m�h(;��i�5�#�@wz-tk)��)Ҋ��V��m�I�s�i��bF�;;���3R������f���d[|fd���uQ�/׏{Rr{��s����5T��@'����ͧ]/߷�.XGc��� �쌽�ɉ�W�� �X�5�c�(O���J�3V�	:j�P.*A���
?���kW��ӝn�D�l$F�-��A�t��}�뛹KzO���b�ּ�!��Y�P�*��� a{Q�K.����!���L?$���!w�a_��u߅�{�r@ �>7^���~5i���=�'� ��
�2�{2�(K�#2,��]���aQ&Z%&�WF����p���\���Z+���T��8'�9ey���:�8�#a��e��*"��!H�^��tx��M��?R'u�ۗ�+	/^�����T�+l��UYb�$�9������]��x ֗��0(V�Q'�2:�_�IG4��
GOmrk�}��eF����l����˹�&�����M�c�g�t���[7��{�mV+���У@.v�e>?H�Dz@=B>G��Adڶ�H*��^��3;V�,��e��pmND�">1;��T���iQ{^SH�:�=QRڵ�z��0�����=R������Z�E�d���J/c���}��KrN�ݤ�$�9�'�5Qn��{�A�xՌB���Ԡ/'v��R>[~Ij5gM�G.�ܖ�/VU�0��t��8��ƶ���@:�y�hg<����{�ؚ#�`֤��6��9��,F�����g�D�eS⣩(y�
ͪ�{S��#Rh�hZ��<D�Z!���n:�q"�|u_�Ԉ`�tJ"��P[���U�xr��>M|>@�ǳGW�K���#���Q��ͮ�
��y���}�u5����աB$F�uSp�ݨ��Vkۀ�EZtqi,���~��{ހ.�I`�����C;��L��"�_��*�}�f�ѱ����M̍2�p'BC�-J���%�3����(je	'� ��l�M���ĶH��ź��'i�٘��������<6_[�66�%X�h|O�.11���F�
�}�Ǝ���_S��:o=аx��0��S���sn/S5��Q5w.�~�6�a0��{�r�g�;U/���yZ�h�9���{w�M���A�)/S(Ȁ|�v^%�-㭚M��+��ʗu�9z�0��Z�#��q��$��ܺL��8�߻%y��ж�����F�ׄ/�,'t��������\}�\ލ��ԬׄQdF�B�:bŎ[ \:�	��t�CU��`�}y��#@�J0��w�/F@H��^�ᩉ=:Q������:�A�A9~Ë4�E��簤���W��z��M�	�/��.�/L�>��np�G������Oܡ�%�H�@���8������h;`WK_�$c79cUz!~��	�̐RI��mY#��n���3d���2C�E��>�d�w�`B&�,�@L�Q�1���>ɨL3�OQ�𷜰��|QF/��j�T�\����;�i��+x�*�z��$5l}�l@'����2 3a�d5T�L?�2@M��Bx����_��2z��6�K,z�Z�����aIx�<��

��O������4'F�ѱ�K�����
�^��P���A�qi����k����O�ۃx��1D�~ ����i#�=)@��5n��1��=�Is���b�/[�@�{Xc��ڒ�X�N�[A&��a�=Rb��D�436���L���wbU4��3����]V�J)�g_�5$��A�J��;��>���;y��j]z(���������.[��XW^���O�h��뼳¯�l`�aG�)ZB`�5��g�mg�lwvކ���/�Cw���P}O�cج˻�Y@9����)�!F�4������I�W�YF}�VB"L�D��~�b$$��1HoG���MA�F�n$��FσVFaؕ=��H���,Ig�-��ե��H0�[F��߷S3%@'�[���?2Q.h_�̓�H
��s2�N��@����7���)ҒP>7�Itr�m��&f�蔲�>�����fy�_[�-G��V	}��?Q�w�
�w�%����Y0ЈP��V�
 ���f�|F���,���6��N��@��	����"'� �+�`���XK�1�h�Q!7����Q\D�sUr������a/���C��qOt ꆴ�	9CԸq��I�)�s�C��Hɫ�����1�Ʃ����7�����,����mɻ��7����m���e�n/�>PX�"Pӏ���mx�s%m'��e:����
��u�Q?�3�h���.
l� ����X��8���O�F��B�G�?�D>+�Ʈ(�HǓc|�1�c0ԏ������dqqn�{R氷�ٛ�mn���և��@�8��è%¢0lLP#�C���:��	9<f���l5�}*ж�E�s
�8�pB�tis����Oy���s�'��!ѵ�/-���CT5 $��W�0���YZ�MI�ݻ�h��(L��zm��+R�����_�� ;A7۾�9�����������R��ᆑʤ��B!�䪙��c��O��;�o�w�D��X
7�5�hESt��h���k-�(jM�_�+e)��7�����*yչ{���PIg������ƚ�M=�����*QP�P�=�efMl"�(�T�k�^���X���h֝��>�4 ��v�}bz#�T�
��(�=Q�saδ9_b�IՎ��i6�����M~ָ�*�Jc��`�������>����ƥ�8��zQ�n�ݼPh3���� B̞$��.SN�,�l�jL9O��F뽞W��F���jdдv�o&e�bcz��:��P|�j�G��T8[�Z)�G_�G��	`�jSi����BN���o�����?Ø�&��x���٬=��T��"��<碞�ND�rL���ZY���qÙ���.�y↶��"���)V�lv�Xxz|�Ўh�J��aG\tU�3��'�+挴9;Pp��"q̀�`y��	����.����>���$#䶟2~�:��2fNw)ۂw��6=�R�'��Fb!X'([bz *d6Kt�*�d vx���?^�P_W�A�ߢ�j9���A���wB�p�lx�%�����eN��"�n�V�KƠ.a��W&���]x���ʤ �4��R4��ͫ[���[���ϩ>}6�S!�6��gvՂV���t�J�@7�j	�M�ꋃ�Ҫ!�*�����^9�4j ���z1�$]va�k�ػ�G#Z�|3P��:M���wN�m��;@��'�pb4�H�UT*׈C-ֵl�Y�3�I�z�l=��q���[S��l��FC����I�Ēz�gȫ��%/ m�V[Z|�H�ڷ���?�P#r��7���%��(#��^�B��eUe$��<� �x���"1q��?�:2R=2͒��	�/%#(DVQwW�Z>2x;N��}���#�W�n��P��Dk>EH0X����c��a��Uz[G*�U�f�"�;_�ַ��}�`�������C޽��O����vcb��}�@G�1B=�A�`��X�J�FK��#�I�F�p���̐wQ&h�K�e���d�X��ڲo����)�<��L>k���_�킞)��S�FM$
뱲�r��Q �%�U�O�����|��]��{V��O�T[��EΒܦ�6�n�W#_WP[iV"�(ci ��Q4��L�r��(�y��/w-Կ���c�z��d)wȲ�x��8�Py��M@�H���&Q�����)�߶$�H0��)@����?���Hʕ�=� ��)��g"������4����P�6�9�e���Ĭ%~��k�a�"���ϦEiA����6Uk�A-��6�\.������Q�Ѻ�����W{��^k;��KxgM���!-�әE��6S�W<8���'�yk%ڍ�X֓6�E�ُ}�>�N�y�
����Xا.q��ʊ���\.���/��O�Ѧ#zZ�����}���~��/pHU�*�ȳ��O��?�ܨ0>1S{o3�������V~��g�FpO@%�+��C�#�k4��s ?pG����9�ЏV�3�W"ކ��cS+�I�qs8z�We`����.�͘J�9��iFZ��6\p�a��du�
i xk�ĀNl����F�w�?��uǎy�*ڊ�̵.��z������p��`c�g�b	g�����,��2��tU�沰%A8�de�n�1�mD�ٲ�腻�:�(�}{c�p!��p����S�V�I��r�"��1W ��A�24߇�ݵ<�OS�-���r��ܺ�iΤ��\�e�^3��Ab��5<-Տ���,��"Q������f<�s{��)��0���(.�Ʒ�����y��� M���$��V��
��e��������^�-[+.��\���d��WA�ytżF���X*��Z$��?���KE��q���ҋe�c�"]e�z�.��2L�TЎ�t�	��e���TH�f��lr��]����g����^��47�I����u�*c�<�	��ؙ�afϡb��{���A�H��>F����Q}	��iq������>fVs�=���fi{L�w��T��{�u�����k_E�c%iT� �C�+*RL>�
mm�}��r]��D��!�M���e˲9��5�'(Qef!�h��X½�����`��]�Q�a ��e-J�|Dt;U���m%Mj�V��*e����Y���~e�S���Rź2�˩%��RФ��	���7�������R���Q��i�.��W�*g���x:��c��lZ�Hv~M�l[^���������;�����h��sI�LX�/Yz�����*�[�7����A{�E�X�J]x�}��]�J`����S�/����^�BrC�~JiTo���I$9�U���"J4����[�ǽh���ĊyPUO
�1Bʬ�[��RU���fb����ft>��i�sBLj?8(_��_��7��Y|O���H#�c.���/�/�23ص�vs�)�Ay���U�����J��(�1��q�^;F͋[̄l�aH�%SW��QK�Q:�N_]����S�vg�mMg����hI�� 6U��'PS�K~~�GTעP-4���<�a��h�f: �&v�s�x��vl7K9�̺�
i�R{J�d��1ҫr�*)�~k��d��8I��sU��i��#����	��r���?|n���hM��̞[�mr�O�?������u=���U����n��=�Eװ� (�M�OS�@�H�d�����"��S���g���N\q@�y��_�2�X��R�ֺw�y�6�0����׀zp�spU�r]���W�i��(Sk�����`4�i���<�����p��r��ƶ�㽑$Ye��NA��
���>t�'O-���r
_�{^���迱��J����Y6F>�EɎR���9=4�)w5D��e����p���q��]#��ȸ��+�	!�G�䭮����0}�Ƶ���{D_��t<dFFQTO\XT��%O `_�5�˂��=}&-��??q��bnE�1���cߩk��8h'�pp���˸b�]� �%K����f��0� �:O�s>ćlu��)fH	YL��0�Z�EA՗�'�`� ̷������y����o𨙁�	{��w�w�dX �˪�֘���|?��\z	�`�����dr�5��Κ������}�����'b[��6��|R�D�<�l҆��;�.l���(nw�j��W8)~3�x�s>��UqA���:s�}}��� b��?�>�Z��=���� ��Us��m�SO黰�eu��h���׼)���@r�bAp�[ҩ�N)����<{؜毰Op�Zj���h���C�VX3�n'*�	{6k�\Ym)��>�ŷ���@���7�y��Iӳ��5�V	�'^��;٥o&�z�cF�[/ '��!�����:�IY˃��,@7���jA�**��G_�c�XÝ_�*�i��|"��&�TۄqT$�������A�K���kʵ5+{�.���:��6��gZ�V\P/��<�+��	����kY*����J��tY��]�F�xY-�p����ӡ |$b�/�!�v�0�X�*�l9��h��_;�<`�f���A�F�Î��{�l�}u����ALNTY�K%>\BX��	�����6�F�|Ù�dL)j��S�s�5�>Hv;�+w�	"i����p��T�z��.�}�1�s�kp�5o��ch�a�q��g�������?��J����v��!<;��X����;����!Y���%��u�\8*#O#;�:��}كL��'��uG�U(Y���;�0�)�������f���*���"�[��n��"��Z�8��.���d�b�`�ګ�n�a��],{³�k���H�6﯁�e��?FY��O5���Ó�,�:*��3wm��xI�P�
G"�h��]W@�N	���[B'�ù�d�yy�	�ONm�*��ӂMd��L���0/��601l����6U�<Y{R�G��~u����#�066�\�����|D�<�2V��(�� �"�ct1ý��~01��h���)�*m���\��Ǜ'!��C����|�˧;��a�xTX�.�aA2�n��_[Z��_��e-�vÁ?5��"~*�l4��No���m�5_s��_D烢ؙ=A.n���pP�� �t�源�k�W~�M��g�����GN O�)��R��(���*�eKA�]�a�[&�xc."\���w�$�ۆ�w���M%s> WA$+��ǳ7P�v�J�t{1I�U���e�+&|�H�>?0V(!��/�\����lQ�zR�"���`�4�7�q�3��;�2�X\�4���y���4a�n}2�՚dm�ٓ�*vΫ(c
���G�Tz�J���w�'�8LP~|1(�O���{���_g�PbFIM���ۤ��E�N�En3V�3�z�J��e:@]�}sN�����D<�Q��  O��~P�ϊ�����J�������?M�n��*#�JH��T0sS��Q�즊�Κn��� w���3ª�����+$��WSwI_�8u���X=�f�d??��d��g&~��D�����È\��=5��1��$�[~Jǅ����8��䏞,ԏk[�q��3=H�نr{.XyAV�	��\VF�47g�:���:�r�������Ks����.N
)Mro/�S��9���)���R�=�����K2`@�>�݊�cƖ!�Ά�-��.��r�tDδ�n6��s��y�d�RH�ݣ��Vw1�Ŕ��������@���=� ��,�Re`;~��>̼+��/�
aF���wg�w�o���yoR�;����c�s�'L��bl-_��e�m�k�uCI~d(��~���+�3g��^t�O���jD�N+�䅐����5/�N���q�{k����+��ΞZ�V��H����Ǎb��s�p%���u�W��+_�l{y@�2- s�JV[�ʢVE���0�<o6�Y�����C�(~���¢�L>TS�-��G:}��6��|�Hզ;��0\^s����r@H����-��A@d��Fˌʞ>�Ow�k,���=�J�g�Hq��8x�7�~}������Mx�Ăj�&9��F�&l��������9Gz�9ƣ�_�# �c�9/��]�G5:����!�E _��^i��~�}�ˤ��<�ޠEBD�^��3��cbW�6�k��q��������=iH[���Djǫ.A�|�o�節��;�j�^`5!�RE3�{}*n�Ǉ���Z"d𶶃�[q�@ȑ'~�PHT��U�L������1�$�l�9`�B�b2�)6x���4�8�M��è{䯔8��̓:��:�X\7��Vޤ:�0��t�2�"��=�V�^�x����l>���7]�C�T�e���[�]�LSOk�%k�48�����$�?0����p�xILŹAO��k">��q[�A�/+
#;C�"8/ҙ�_��0�[>���Ʋ҆ԉz�0o�/����3z .�!��-*^�k�6pp��K�����ī�h��
rM�����1mc�����ڍ�/�s�j�f	Qc�g�l>YGd��L@�Q[o�g�pD!H�0�X�G�?�7~�-�Ṛaq�^R��
K(.1����AK���*��X�o��ä����5���k?��,�
��M���ViP��� S�Ov4��IS���f��'�eT7����!L�1q8�u4��<��D��Ap�}�����)��	�J�~x��v+��v�o����?�b;[���2��O:aeB�o���q�iж{>9��.T�r�q����t	����t�BKQ-��䂞ʹA���f�ӈ]M�I2�0��<����~�C��W�2��ժ+�G8�$��� ��7���D�\�{-�c\�O��:v!_���S�sP�+ak�HL����-<ɓ�n
��HR�a~P*%�#�y�u�pI�H���ï8!y����|]��@'N���i$W������R��2*0������+b5�L��f�$�`�2�1����s�APJ��	�a��%}�托,}@�.�C���lf2��F�����V��Q�-]d��Ӧ��j"���\�Eբ�1
�Q�����N�9}g���+�o���J���� '�^R�pQ}�έ0��.b�O�m�Gt���N��̷0�W��C��&������0�J:B�"�����'ܒ:�j��cEYc[Wn�8��s�#\>sO"�����[� ��RF=�����}����/�AI�3!5k�8���u��c�i8�U�ܔcl�_WӦ�{�𩺤��e"	RXХ!;�RߋVU\�?OI$��3��P�|q�L_��^�2i�Ù��A\!��(:�ݚi�c�"`�88b|*b�p�k�N$6�hW�-� A�B&�����T �d�=m�Q��������Q�-V� U���?��L:��!���v_Zά$6wZ�qr^��B���5�ۋϋ�������Roޛ���&�VS3��#�/��?U[5���;�V�C����BRIO#���A[��״W<v�Q��8W�sl2wR�`�jȁ�y�U<�kDf�+`����P��rX�G���4��2�^�vr��Gb(���o%��N�E	������͸vqKe�WU�Z	���J��w;�V�_���͊����y�o
_���^HΑ�=e�y��/��d��I9�R�9����l��g3��x��\Q����6B������^�mX�_�5fǭ�U˨>q"maO?<�x�J�70͇���Uv-�hEv�4��[ĒD�k����2/B����#����4�C^CO��\�5f�jR���SɌ�ٯ�";_@	�Z];ٓ������eY+⺳˳�+��%�-[_ )���kL�ߚ7ӌ�#
1�ǅ0���_ph��I@����}"���] �ns[��]=� t��hH��R()�LjK��C���fD �ߙe0�mi2U��@\3h�fs:k)�=�1u6�=��F��.�t<)XKtb���ss D��9�p䏻��[Փ��̷�����	U<����챳J|W�,��9h���IsN�+^?R*��ĳ��M,���t�\U��TrX����+�zy7t��Y|w�S�,=7;1�	S�Y�:���g�G����Kx�B���I�Q�~����NWFL%��"<�9-�/Z�쎴{�Lr>�b�&�ػ�f��/���`=6��K�# ���ELu!�l5�%��v�U����rN�Y�\�@Y��;��3 ��)��g�j�!6��P�ة�uN�e�p�I�&c��c�g@$
��{v�(������s�&^��Y.��`Ƙ������������ǿV#��rP���ږ$uG�h
+�ɀI�D��Z�3��%0�'��A�z0c�<��v�@�ÈwƩ������4���}_&>W'Kg^`��v,���ޔ6�l�*ΩSw�|ٚ�	���żO5�a%�E�H��� EzO��^�E�zW�}MX�qa�UOݛ1G��JG�I�-q���q� ��8pqբ	��/���Ez*�t �|��2��j���&�i�=(c�
�	)n:��N������vA�r�$=_�RG�/�o�a��N��W�	aO>xO���Dt"�	B�+�O��O��s�����XD5>�F��+V}��)(h������T��2��އ�5����D��x�d��{�~�y&��_�I${��\?��"�*S��<���b����鍫H��0�֔�y�Kx�![�p�;m͋��_%֜����Vt�al���q��b�Hqn×(",��@$��n�J&o��fn�k&4)5�Vk�����*"O:��g����hK�Y��d���Ȓ�ܜd"���ɋm[Yr������O���s���v��dn7���	:��P��qDgź[>��ͥ�8H@ %��D��݀��"��AGR��(	��Gz�\vğ�f�U4�/N6� �P�(l௷�p����B�����ݙ��������f��P�����fe�͈�0n��I��]�PhZ�n��V?��@6Af�<�˷��whlի��0�\�s�0?k$����o>�u��e���~nHIE���n�0+��{�k�Q���X���jBg��ֵ�ړ�gT;)&��q�Z;"���d��^�(�"����Nں5+��~W�֠`��u��ֶ=L���ϱpZ^�_4B\���>��48�"e����w(a�=��f�'F���O�gB\n�Y	���X̟��`m^#^���y�!�/��y� ����4'@c�l���Ѡf����p�5ѥ�>4�Pg����S��~Oy�P�0wX� ��E#�e����$�8�սep�+G�'����@�,�w�C`fI�wd/�iCv�	��ڝ�Ǣ8|���_ZI�_�
����u�TIU�964���g���]���.>����yo�~7{�c�n&���	u���=넙/��W�<,C찐ŔqN��FRvT��ᝒ��e��ot�&�Z�	��s�%�&�ս�6<`���&_�>CV�Y�i��*l{]��.�,N���d�`t���]��M� b������}�wd�O�iDO�N�d��ܑg���?;��1(��s{�Ɩ?�m�VK�U�F����J)�6n�b�}��Lĵ,.���ቹ���,�`��M�:�v����='�9����p��+$���X��c��D a���Rq�gYMg����)�guO�]G?���(	���,������ks��]do �r�ތ�����@"��/�yG�xY�o���	��3�7��'{�lI����$GR��j��1"�<���b�P��狏O�4�wu�]l�7h�������k��e���y�Z�{��V^)�2eC5����Ch�gy�T�Ydce�r�<�%���"�ݨ`@��FŸ���Z�u�k�/.2�\o���O,R�3? ZG�"�.��K;"iuT�.�ָ�wm�&���X�DY�B�n���;�߻M|Q�3pk�f�n�}�T���Fvc��8����[�;R?�rc�v�9�%�t|�v�k��&(;}y|D]�9~k���W>䲦9_��ٺ�QێŊ|N(y�c�LA����&��a���_���Y�7|2%�rP�6;���c��)G�{�cw{p����nܚ��Y5#e�b��-�5�m�����ޏ'��|8���2p��97eH[�NP1��k; s��ܜ0�N�m�=�����uv:���F�����	҇_<P���XW�F�pg��Ƙ�vF(��Hn�*�x�\�kJt��"s|v�7��3��5l@7�9i�M���s|̖���:�:���DO8�R��h����Li��w�F�·N�0e(��� ��nӨ������H��h����2�I�x��R�N�枧���k\0�؂�UvfT��|1�4-/J���<z�53QR��Ff��ԫF�洙M/����8,�Mޝ1mJ�yۛ5e�Q"�{{�&�.�H�}����:��q�l�?�_��s'�����w@�[�d�QK���=7��^��PN�nݜk5�u��J���^q2}8z-�8u�4-=#PS�d�'"��`�JE�H�^�s?�HJ3��Zj�#�\����!Y�m|9Ց[�-�Z\0l���`�Ԑӥ�d��q�^IfV���"j���h�h�x��1˽VŬ��?�{�v���+0I�;���^�����Qs�H:3��(I�����շ���@�A+9��E�0�����e�W������C}���(NW�v(�R>m)7���t��7��*���P���Y�Ļ���:�Ν�Q���@����;.�@��,�!�}鿝 ����hs�x[��4�f�5�^a�ؽi�M�G{�_X�]H֚�=Č`U��V�<��1��^�d�׈s���Pv�FAȹS���^��k|�R�N���1?/�!B�51_��ñ�E &�
�'�V����u�S[0ԫ�O>��mkd������j��c���cs��������&�"t�ss�1�����Z-��f�,)b�E�S���w�F��!��"����xx�Ñ�3�s􃿯r;�u��0��ZY�x:3�e� c
��}���_�>_f_p��vr�r���i������F21C����(�:l�}�5�FUuh]T�P��	z�N�br��لɼ$�Y���#����
G��	B'����μFR�̌�_0�����A��
�]H�]���#���ປ�E߻�ݜſ�-&խP]��涤Mfd��P�J��W����a'�V����ä�9����!8�߈�@i�M;�,4mc���Lf;)�;�)e��2`�!�������\�%r��Y|�_MZ�{@�6� r�,w���PID���K�1��9�����e}�H-��Is;��+}�Z1��*)��o4���d��vÖ
�#��p��$RA�(S=��?���N\��YyL�?��v�mn�'/w��~��=%{��8��o�����KJ�::O��5a}v�`k�m�;��2�~/[jy9���e5.FP�Ŭ�%T�=���@{c���{B�1>*�B���'{��峜G�[��4w�����TCF3�k%�@�i:��n`I�P'm`
3G� �+	�&e����u͊e��!󩆚�?��W^�R�
'%=�N�A,����@c-�W&u�M �ojm�Y[���i���L͝�[�Vcb��s	J!��}�^�B~���B}��
��h��X��$t�M�����%Ep�����$��LBN6����͠��T�*��m�3�yuYo���`���.C�rxԒ!l�w�k�8���t�|�S`�{/[�l�DL(�����i��5lb (/w�� ��t�����vS3�����j���R���,o�%��w�u�b�U�C�6Y�7M�e��&���~��vF��ڭ[����;|�ұ�.A�K���,g�������c���m�i��i�����|!���9h��6�|3�dpN�Gf��:�7D��նDC��'����x�q�\�-���#R��?dn��̪���&��Რ�X@fg���j�x]���V�h�	���)����R������]�"
#���?�A</)u*7~"�27�hbZ�x	����H&#�x�$(�&��]B�Ñ6a"X38Ԫ7!˵O
��K����9��<�5�R���/|:Q���Ĕ���@k�1~?�J�gzV�`�XQu��x`�FY̚O��:=�E납��H��㬡D�䩳Z����/���{�z
������P�H��(���O���Q����J4���[�)�o�G~Z»=����	�b3/�~�7ʤ����o�ŵ��Y�N��3Z^�����0b[4�8>]��+������Y��z�r���NiT�IƄ7gu]�P�q�eR��?�S����2���s���s,�$�p�%���9TT�$!~��xa� μzj 9׫)� ��*3�d%���ʉ��!���3p����</� �[��z|��?��cI���=�Ml3Z��
�	�G����s��Ӫ�H�l�s8p�z^�
����D�>�I�t��X�"�R�~b���s�
�=$ؗ�kr����P�TJ*��T�����y8��4�G����Y�MIK�r��z���5�`W��9>9��JZ㔱zMr����Ӑ3� a�ߓ�k>���Ǣ���3�n��D����4YrPol�2��P�S|ʶ�>��ۆ��Y��K�������Vk�3"�9�l���T�.?��l2`��]ܮB,�l��P�=M9�?��9)��r����nI��q_�=���m/{X1�g%�����ڌq��[	,�	]v���$�̈���y!K2���#����K��i�hmP�	�q��jA�Vm�ՅW�L�+���o:"ӥ_�^��m��X9l�kB�p=�8�)jA8 Q2�@��fA�ͫPi�s��='����BDZ����o�"����}s�Jʐy.w/<Y ���q'A#b�`�r��[i줢n�M�g4�ܗ���[�F�˶>�x�!�'�� i|�^�!!9�8=�Gl�u/����#�&���d�s�|����dm�w|�H�v)N��J�����L�*�ոM����`�K,<�S޵9��K�m���v��
8���1-�b��R�;mk�� �CdZ�aX�����/��_�H`YJ3�.��.>#e��w�E�����5� ���_�9r���Ɏ��ʦ�,%�A=��er�S�N��E�ٖ>@8�;�-�.��1�y��0������I�ώ�M��YTi���}�G���O��yy��D^A�ւ���yz�R̈��q�eA��	���=+Hjd�B��-�#4�<a~5�Ҭv������}6�JpKx@��$�ŕԖ�q �aC�qB�fM\��>b����k�~��Q���P��4�R7� k���8̤zS���"�cF��.(����"�cA+���A7�0����_�	�9)���i�E���z�}�N�I�n5�b�Ƃ�pg�|�&�@��R,e�Z���*�pn:����DSyۙFVh�y�.� !�W㋍��c���ݗ��_��t�ij^j�p_j@sa�b`͸�*`��`d�8E��T��ʡY���z��_!��ź���~-����B�Hݶ8%Z[JA�Ż	G��b�]�H[�m��π�Y�0%%5�-���~�C��K�
p�t�߰���9���d��W��ۈcx��:�ԫ�����;���<�ǥO��zB�SJ�$s��]��*"���U�z���;})���	�e񼢷�NcY�;CHCyw��IH�2i��n���+��W����d}$��R�~orC��'f�h�gNx�4=�cG��.9��}T,2<�����*�;5��k�a�u;��;0����O�?�-�ϊ��R�_����h��T�d�
jf��A+�� eUR#$Fkˑ_M'���s=wZ�Z1d��L��?�$Va�J��w���.]ӛP
;��l����uGT���=}�Ë��!l�/r+dQ�J?���!�z�U/��R��.V<�B��g{�(�U;U B� K�,L�p���=R�����TU�&>�YL�r�6�.,s�6�B��L�R�/���Z��s�e��fvr�ղW�T����fe�m�bE�fZy��9���I��WA%<�r4��a��tiD��ܷ�rtn��8x�����U��������+�,��V����(q��/�梬v�/��\��L^<*w�ֆW$Y!�WR�%���<\�a�<�A[E&�P9��Mn�!�
_�
�f:t�( �UX> ��1�)C����c����k:�)��gU�CEf����< �>�V
A���D��o���5��tY|�Y��]?aH�No�eo���*#���@C��h�"�ߧ� ��u5�1�!��1f���dXdܪtK�1W����`m����lk`^�Fr���w�b+R^�h����
�������s�I��������x$_e(B��8]Y�i����G��X]&�ގ���w-�n��Dm���ZK>D�z~3˼s��s��W��~���J=��z��6����_�n��/spL�~n�d��f���j�u��"�bz�
C��4v�ap{�!'u>�U������OUK���hY�����E�d�t�|���J�z�a��uu�`�!Q�k�����l��\G`�Bs�=虨ڛ#z���z0,�1�@Ǻ�N�9.`��-^,�gBw�����Ț�f&�۾�3�r2��h@l�o@��߰So��q�[fQ+�X�y�H$���U{��[7u5�X�dŧo�3� E6M�|�@p�:��$k_�7[��)Q3�H��k&ٖ����Y�V���^U�ym�ө����= �c� �s��v�w�yKf�����4j�<�
�����N��;�2�!�wZ:X��pσ�Ħ
-w�Ԍ�z��w�gÉ�d�
t�;�����=�a?�����"�rr }�����'~��cvs�[���I:��2�a�6l�Q�Tf ��x��=���m�F�^�.��3�&N��ͩ^�B�C�{� =�0n*e,I��|z�;{���%��^�jۻ*�a)��0=�]�O�H�Y����i�.���aP�j��FF�*Ve3X8���<�����='>>��a��j��V��C�C��?��h#oq+��\ �5��g��rZ��.	�w*-��Qx���;Ŗ���6�e6?ѐ�O����m���;��&�DݞRqn�r�&���jM�T�F8F"q��'���.��$��p� ܖ�٦�|-�	Ւ��� �GQ��&�Lh��/�l%�=	?9���5�)H�ӇW�Z��<��������U�C��i�'���1�`��J�ȡ~�/c@g�j9U��L���$�����s|����]������]�Ӧ�e65��h;La�)�S��C���z�����0E��R�YW�>lfX[�Y7������j8��R�4ͽ���u�W]&�fjK{`���UdK��X�b�svU-R����N�B�>z�.�ߨȊ���I�;����PO�z@ ���@s����.�;�ɈY������Y&�N���R�,|x�_�����%J�g�AB��\|��r�/�F�>�IhN*,�4lX�וJh�)�b��W��x���=?Y&�(F~�e_}��>��^ݜD5�q��B��G+L���"_��t��������%�کA�ܦQ}�<���s��懶`�M2J|�^� Z�l���� ��8k)���`���)���sJ;��ͼ����Z��������.T(�&EZ9EO��@��Gq������68��x$��g��uo4�%��ڶ�)��P�-z̾`1����1`��>u��Y{��p|���K@��#F�2[�ۛ2y��'/�Iv��.S��l���GԊ��.d`r��ڣ��h����N�M�<�/���\����膝*������{��iہ�_>qy[
���Ñ�v�V���c2�	DO\?�U<L2g�\��ܼ]���+�Nu����