��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊"3iP~bE,�ﱃC�1)�/f5^nXQ3kP�;�B�xi��+*l�/�,G����(���)���1n��1Rq7����� �i	M��=�����Va��YwN�"(����N�mEa�����x�8̅Mu�w�����RH���f������D�b�~5��>
/��$�(�5,A�6&::���w�#��`�^wZ���H�+$&�{k�W؍��dal>��m wXF���ԄL쑩��л�dR��I�&1\�Q�oI�U���\�%2�1��s���h;k(�z�c$ y��
,wXjz�̺3�BrN�a㰸\?o�3v�iVQ�y$G�&t=���2�g���v�N���.��oyw��
m*nf+�h���ñ�1T���-s��>M���h�3�y2d�E�j��[z�ޡ)P��$�w���̭�K�F�w*b��oZ������w����l�s�,�����Y/�@�aՉ��t}X},��)�Ԓ���,�)/��������kZ�}0����̎����D5���Z��p؁����=����n��v�����`6�Gپ��i԰��#�+k�;"^����+���:��_��\�G�k��'��!|��Ч��侶T9�_D
�;A�u��i�8�sl�5�O��P�v U�cl����N$�'t'!�N���;�~3���r�����>2����XR�i���O�IJ<z��gD�] W;BUr������/�hӛt#�rt4�+1H"g*��o�1�	CSU��\�.Fx��� y�W�ܼ8��V��+����fuF�Č�. pnJG��`Ud�m���+Dl���čP.B==�``ri��T��]�	u˼	�dŋ|`J3	��!$����$:�Y���192g�;I����ZG@�c�OC�^��6�!�Y���p3{�,(~�����w���������b�>�)�*U?��� 8�Ή�\
S��q���HGV��o��I��XC�l?���23��I�Ւ���]�&IunW%�9�]��SR��be1΢��aK��-�Y���l�X�|l���]�2���3[r�*se���|��b�?�	zh���^O/�<��-�����kK�$E�I^��!%(kC��O����&�A_#k��WN*j���\cOKD۱���Ag��*�,2t#S;�nW�t�$�d�o�Z�Ep��*�Z��~���d�u	}�-���-�?S� ��o�FR���B�9�,9#�ƒ���g�d�4��Ѷ����u�����L���Y���2#���ѩZ���(��ô��1�
��j�j�ޢh�m������")�O(�������Ñ~+��o	>ǒBJJ#"[��N�~�T��9''�Es��� �G�&���-ZY��tQ�E� ��Ѱ����f�v�9��K��l�c頕M�JV)�9L��P�Y��.�}
0ȀQ�˕%Y.��ї��m��|79��E��&�ܫ�9RթR�Cع����%k�W�_3�M �W[]��1[�u�>`}kϵ�\1_[�{`M����T��^	�L#�Z ��ڥTu��æs�Oo�|޶�-��݉͞�E�<�\����EC϶k�X5�J�ޅ�B�Q���a+�LPF��`����笒����w>��(��u�{sx�q����м�G\���Q(�3�_2x'F��J�0����-�&W�M���� �U �5m
]�@�+B�K�6�������<�a���hh|Y[G� 5U4j�z���ۥ�Q�O˗�I����<?Ũ��+�e��di�E��fzw��jє���j�sS��L�=4�㍻&�%��XwF%o�?0�wJY��ê ^�hg����L����talZN��`��jYk�lN�����T�@t�Nl�N���`��5Q�H�`c
c�#��$�+��Fߟ��F+�\�q�&D��c�-k�ꮹ�=�>��7(�?����4m
Zڷ���e]��0�d�VF�׎�$�J4�q�)Tޣ��ױ%���,i��)�hX4{��lC��7�	���Wud�ΆI(L�L�t�{�[�,�O;�b �Φ��"3Wf�뀚�C�B/.� �mе;|w���˷���j�HV5��d,Il�����	6���u�W���ˈE���Қ����&�PP*
�EP,[����x���@mc�[�/Y�"$m�E��3N4X��+��ޒXY�á��6��.V����g��A��Բ6Df�8��>�>��iC�����>9�\�ڈ*A�]�ř�?�^{[�LbP����ҋ͒Y^<R�n��ܠ���7�1iJ'Λ徱Z�3=���������[Jđշ1�� |Q��XD��t�L°M�<"���ԑ?���|pSqǊ����|�{�Ձ��3�y�� ��� V1�(
�Ԟ���U�����m�~�R����A�;Mv��1�e�����b�'_A�\��bD�Z��L#�7�3�C0�j��s��]���SS���	4s�PϡE-M���K0_����W;�lČ�����x\�S��v�v"˽`Kh�&2��)�V�sH�`���O5��N�!��h��g:�`m&�[B��>�Ĺ�=*�����R���?�!v��]ǺM._o.�Ԅo"?�'�su:��_�}�)ߧ ������k��K߆rc���'��6Q�,�͡��s)�qt��+n���5���I��`K|����W�)~+���9*���"K��zZ�Ȏ����-���8�{n��w�	�/��Zo@� �nA�@s��		6z�|c1X���Uwi�s�ր��(�a���j���h����G��7�1���0#���w`qxZ��8j-~O�D�z�RQ��T����Dw�_���[��G�<�#r�X�QQ���W���5)۽�ey�i�j�c�,H��g�$����X���R�L��>ɂ�aҙxc�������8@�9�rX�zD�U������/�:�vɯ�Ѩ�y� �8"]�@:���k�dA����.������ ��i�����4��[���p�[��,B�~�6������ρ�g"Y�`<�W���_��.�֬a�X(�z�]���c1