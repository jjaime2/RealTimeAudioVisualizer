-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SIClsRQEZmiXFMJCoE/zj5wrxqMrVhKDHOKeXciOzjwKczQ4DhvDPdXhJ2wySv2vXHUhhepvqEGC
oWNGQqHEWJ0x1K1is43U4lt675Dw27lDN3JX//aApXO4AsQVXqPMDNtFdqs1eE4kVJxfJ82EYDZ3
UedDjVe9IS7fFBdaIFRGZD8racEMUP9y+gEapO9/b2qLJXbC6O8Cll037jxqxWFKs6RJ490XbqzV
FjssrTLIlBXlOp7GvcxUcuYU9fTlYe4Wev+Ztqh7Kyej9rj04Q2xEvmA5aYWlQVR9lNrXiC4sN9v
cDe0p5jYcfVRt4OTu+imQu848OA1OmoaI9MusA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4384)
`protect data_block
uEMnBzdatQthdWOkYry5TYjsA/UgWRnXHKpbH14U6DbmdBjig6onqNI3k9oV7J2sPHUPXGOjqJqy
2PbAA6TRzucsuMzjaHAw4mO2rpSbGPUd7IJZnmnnWWnS0aw4+SuxKs+ZKtfoUmxBZJ3FfIb0KTs5
RyVJt3YEJdnFGDqLfUFMP8EUrQdMbGnA8MsNgBfuN2xJK5HgRbHcHSiZ2R/5s/1oJEwajHUkgSU0
ADXaNR4KJTkqjPVsmaIneH1QNVGK8Hjh9KmOU87NvEMfeuYIe3g3x1D2DDwgOJNMlRM7lm8DiW0T
WH4tch8beFxBkNiRNTOa4GxgwHqQSqajZjWt5PZg+ujV2bmqlffqYyaMo+5lrevenJnYaq+1Mrv9
PLGSnmQh20KFdgG3gXSyLaWQTJZQm2QFQ/3k5XYryg2FdGGujJcBGuQu9uBAcp7uphwmGOAJwvLK
u3nhkPfTTW72egK5CN8xoB0Z60vQJqVM7yAqMvaGgtXBq0bG69uY3eLrOlUPViWhEo8xKal1v05x
8m/5utPv4cL7xw2hL+eNDdigkCQs70X7OD1KrDHpRgiZ3oioDnBpYcIu6BMrer/mDmLPTn3J/kgG
jMU1qm/MvBs0mPeEp/XtfUFwfrDODdfXvcL1RIyDjYZ/aT9DZf19/SWu92LboyayXmmFKGDJdtdP
oYKod2gtCkJ3zSNao+3XTaLCu9sCvbS/aqSwSmVHTUmE/OIZix0jOPwVqjcT0OQfcy7Rjav6XVAa
odad3y+Y2ckMZ4Zael39JvBLnu1mPsoHH1kuNgCTFPm/uzThGVFbDya2B7Aiaj/l7msqUKb5ZXFD
UNQOKlkR1PJ+pvSP5I5g7ka0w/LC0qgTU2TBQcXI7t0P6EMMArPQDvmPHpj+ZA3H6sNKyt727Rd2
Cp+DipWvUmYRcxPfoGP4xRgqjl4ey76NblMsQFRkEuN4rCApZB3SwaR/ExSJAOXyarsjD5HT5Sfz
4Hu3XxS+g8jKHwOCD1Jr++oXy1US2q9fjYcpNUkfX2TaBrJ/Cl+OCWE5U80TJJg2B55yQeN8Fti0
zIiaSZhgYt7v+x/5zcbjaT2b3xYFDK9kmu/QxQtN0kNZw2ceOoIay0gaKDZ5MAorGfCV+/5TTxBy
7tE8TYq1pfHduv1lPSOtmLjLhbcqUx/Qdl9Lo9l1FGSDcNBW3pw8OMcPLtTHZpe312sj6kMz3QcN
/yMXf5A0M9pg1qiL0Hjb1xkr1TTATekbpAI2nvcKQ+j3RfUecdCsmvxcXQk6pzDp5XSQoUHJgZhe
y44cRPvLDGUAJLnItu2oC4OmuyPXCDJp8Eo3B5MiXtKyRt/l8t3q4AR9P6djGsG6wyBzICHHOJ1+
EwT/T4ssRl5uPdZ4/CtVkDKgK/YIcswmXlTXpA6CTJZa3hWKrOPGcpRXuYxqU+0icPvPO7oR2tBq
745wunt51ZEcADtnvQYB4A6XV5wPjv5cLtX8eRw/X0StRoIcPSiBCqN1kVh5L0Ehrb2uP5rpSRg9
EEMOAUqvIoa+3EEW1rXBRknPczcmEAxn51XKyxvUQOz76N1620WwsmNQEKJcA73GJI38akN9Sfsi
imWMh20cZ4c6aYCNbeOLcHGziUulAqr1Ma2nWT5OZqnZuPor73kDBUd5DthBZZI+8afxSXKDNtb4
I2AWe8ekHFcPYtQH84UIHkg2GvSaswNp6OOAcbUYvSosywuWxxpXAYGR4jZji+GxkB/czwaCiomU
n4ZyTVJVaD3MI+NxBVDyWfBiGayQPC0RS3BvbwavJkiKDmVDH3ZhWcjrQVRA459MsNWgR6TBiZ3g
6ApJIb5MPlgrpB23ATvzso3xkudFBJA0U6MThBiMwhCyHvCJ+S3tU+WXg6ydDM3/W/mVl3cthnuI
ktxlIZzWFeA6ndJkPiSye/Y1AJnIDi/2zVONAxLpaOa5S60t1Qcx+bzXHCTDkzZojAPTZEIxjZVs
KyQvyfvXW9tQMFDU2x11soUlY1CwuGZHJjC0ivD+9FuZ6w7e2k1lwdZwy/alikaxAyZ47KH+cVKe
jdQUbWDrNx5J5VbZGBfaX9csX0SGnO5MsO5X2Qn6R9DhigDdJj/P+KVpBLSgUjH9lhAVBhab3Oet
jsuksK8XsPrnRm3a7BSouqqrTZpjeu6R70iMne+7+XEMP88TuoWMNVRPLvbeDtzNlw3bGjcClVPx
POqWaM4hA+gwk8DZrSRGoE0uk+G/GPsxmg29wNtwpzXN1sB00kPbsUijyiKiX1yEfuC1D3qe77ef
/YSwKevb5Wtbu0/SFmNZax14SMJXXd1MDFan6C9GihfHRledtxctKIE2shn8+CC3Tqqc6IgqQQhQ
YWqyrTrmIO0ExK6C7zrQM4KdRw9itYmi32GimaPexmd17NQN0NDrDW8TcjzuFRAdSDo4Jrb+96Dw
JRFt/8YLGTkIYlRUgsO++aaJhbekHSqKp8FRvyXs48X702RIfXIEAiky9jxmSAGX8pSeizQBvpvA
DY7OtLEqMYtrc4/w0SQATXWBankW8z9TXdDmZYzGBoZhniVcpJMscB/pf9DgikBlhlFWFkX/SsFO
m7xDlrGR1GnbAfnbjhbDaIwnGQ2ZQwCf9+MAdD33XgMjnDl3cVECI0EvoXgtYV5svDth0dcKH4M4
nLAK76Gf2L7pGNGsWdqG/k4XRtHcr5RzAVaSEGnAObHSXc29iL9Ml0GvOmGGPkQ+FNeCwjcsbsnO
wLZjTT4B4YjWFS75VEbjwK994U0kJKxx8rdhslidS3WosHJyVirJklUcr9pDJtSSoO1RKRHDzKs+
kWyPg55+STVJQrW5JmW1YShGRGQWA5oQZUpiFgzYgFu+VTCrj+HiMiDsrENseibu+/ACcNO6Mx07
4s7i3x1nYxVLOTKZZZHTUK68E4S6NltcYLzh0zqq9Suy21VWKi6C5n7t8gpA9+r6q23B+40noO2e
Fsw+dIIvb5kUKFaHDVw6uqdwVrjG3lcw5RDnmmZa42ILzRhI0Go8jDv8bL7lzilfFK3XtlCbsI4Q
57Z4nfKITP7OmK/xt9oAWz5VHFR+ZFOiCTCZ9+0A8HdLZBfYFlzoa2MvkmssXE2KYpzxUC1tn9ga
be9inr5UeXMG5xCGf1ozi+sVXn0vne3zuGg1pXj43Ai+rj0izupGAn+sgensaCAuBUtynK+3l1Kx
zIGF+n6Gj5oitBtqmTqW2zzufd9OnwdX42/QP6+YD69grjez82ZyAMwXVSdrVRn4twjfLqmTm1Ty
CxokGKnM47h5NQEgpsMLAuqYTmb2Oj1Eo6wxoXRtrFyoIyb+/2RCtjxewqSSPTkySlsOEj+ZlmJx
zH0yME9xhZtt3DCO9RVpINxt3yVVdPRstk/QOwoC7RQCsNxE6l05fGFXqU32khHV5jUxQ+sZUt18
dxwzYnciMNyBW6u2/wg6Wi2M3/RD8wMlSwTryqJuwM/dpgiYKaw+9vQb9Zpe5dh1TeFUk31kiMUL
iMyuE6j5P0d81KyNv6+rv3G7dGc8SDvucV+VjBGB8uDPy3NX5keNe3BtZU3ckQdc3LSO5aHYmfsX
T94OOPM52kvX/iDqKwOh947gcU84yntj+XdzhULtOUS7jZvZUem01aO1seSA+6nEfDv3wX0VHw1E
zitJBwYaLHywOiydxwSyHMdQNuWpJZ4op48dUire/vNtTdMmmVIXi0Jpe9msH/NPIvCQQXLHLLEp
aQdcfIZ8DFkfdT5la+IO5YWFAjYgSXY9qVj4f6WnwJ8VurCQ+DlEA25SVq0Cjg+jvWA92rfkhRbw
hCSVnjyy7fRJu13FfvH8eG1l3ldHYOsdtavwo2/9BON92e63b2HkdXDO9lNZ+LREy1LDcxMQUcD+
zBrx9+8o5XBAytEc24QvFdlsM1i+lcN81TCrZ0J1TX7adpDkUcISHwyZFLTb0scnm+4Dgv/OoKdq
hyowbIiBg9CEkzRooEtsIq/XAGgu6r+S7ABPjcwqmBWjeUNGkFPxtasRod+fSYCaapbP0g56xnVo
2K8yraJA2F8EtJsZm0twa1bJpLXoisrvasttVLzM01e1R/zH/h6I4WgouMGHzXzqTyGDlmxRx2hy
CM9CIKE80RwavU15red3rCZjbOwe7Ub+DTwDgV1EMpTBJqnH4PfRCQJs5pGFG04sRL4ngJ2H7gGA
QbOApdHrLV/1CcKaCj6TN60vVv/4iJgkl8RFBzBR+QlT8DPJ+k9dsnBERz+tzKaaQFHunugHYGXi
5hogGz70gsAHPmGWP/AnL2dZnGMPva+Hi+dVuzoqARn49BDO+YSKGm/Hga1Aq1wJ/JqSqZtXjXBR
Wwf1Jkwad1cI5+Ru+EjmrPrnuDSxYWzUXKgaybzSZybYmTj9w0V3K91rjGCI7afy+dlbMa7Ig7IN
G0zcWwY8K8AtiHDEzATKSVwF1ajCcDwb+SPDaI5udAbVh/VqfW9C7KSgwuuFhqYm2QRqw2u6k6Lx
aeW/2eF028Z98pag3X7LvNNVaGYCE85fggM6PWRaF+Bt9JPOPPcyri/538s21p7OZm5nxAY+EZBU
JCkNy06dDXpjudbM4G+lK0HPSw/D+xCFcATHHp5/+SlsbME0Cg55HcemiR3S+DEwaG/+chgEnnt5
wsce3P5swuFUSH6uBoHxz196avXlW7CDgy3sxHup1vaMx2UvcvbZsk7QbzhY2TKWZkgLzjl8aRHi
Sri+cAJGdJad8KrjIBTdEXHymOoP6b5yd7zHsXvVDWP1aC9Z1o6AddQPEk3Vx7sewRGkJl3hDsPY
qPCTLIBUWvt7/GeGC4mtqGFscYM0pxhUqYlH8MAbdMVVznfIiHxll5cPQMvMIt0i0MxreWkSqqSf
cMI1fnJkjj1CL2OVS2Ng0o/JL+xWrScKw6LFF/9taIAi92dcHGlKYkV2EslpAudicMce0mUsTid8
NFjTz5FzmE2ZNU31IEeM+LT4CU0Vn38XDmzCM99Asm4yjHpMnqtI2cgzvxEntTaV7rpQgFbM3fa7
6lxmyJMRxHrC4U/ht3qW/+qNRPyEHd0OeHqh347fwnXiSMORDNVQZ4d9MapXuF9liXlv6+0JeLlW
xFMZ1aXIUozPa9QOPJa0TS8UrhFGF5g9c8zvVMYNKL/txfUTbPhtJn3yMpAZ8X5B9VdVLfsiKTNw
gxc9B+N9LRO9FnCiSSZm0Z2OGGZFwuIxNkLNurSWUHdm32Qtb6xGx07VZ+rGkpBklR/8pgZZIuIT
nQQyObAa+kj+4e5g3bD2mwtA4zUaoIXM0GkOWh/+lmg9Sf23//bmDlTEgcLuws1WlVrSBA+mL70p
Fg2JCppC7QXMEnKtHyUscI8qbPXCyry/Z3q1HEl7GucCXKR8QJt1m128OgZ5LpBp7laozAwW/sqA
CjhF+MEOfFkGac66vvA+mSYuAG0jIStu6s0gGIh9dSK7zPaxGXL3fzZxFCHxHdH2QGw0lcrzz34i
cS1dNlZyClJu9mrncHgrtuWyJL9r/OqXat+RvjhZcQ3JW1GGGOXl8bZcEDTwOCWBIZH1FPj6gRFH
L0AOAfCaG7lDwj98cI5gDOcb7rbbTxH9v3JJvTBYVTKAJcuzrFq3N3yLr+JeVk8UD+i2xM17fPEd
yG37qj59f6dXRiyiuWLt1J5xWN6i7YoUzRCndi973L+soCHuyemFWL3RTyBBdGeKDH36Xd9HxmOb
pW8ubL50UAGo75a8tJAqDiaThkn3cb/Rv8Z/fV/HJEMDnZU2CkF8kVcOs8tVHUyjvrERgFk0mZpc
zsZBkrA/cua7Jyk4a7DmcrLBs5fT1lYqWm/z6se4zvokf7rOcvV4U43Mwc4/07al9S8QCg==
`protect end_protected
