��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ���l�$�'�Z���u��E�a ��B'v/�γݩ%5=F�7z�N?ysV�k�b#!sI[-~�G�m��]v��G��&��qx���m/�H�w��V����f�Զ�vp��B��\6�Ads�-����jfc`�kQ:�k�ɭ�|��&Υ�B��n�R3l=���]�_���Ro���*s0��|Ft�m
D�e4,�t�N.��a�˽�T'�C<`�e����E(�!$r�)��}�����3j3Rċ����7@�(��zmt)�`��L���Ì���j�LWS�g�K=.���F�-J����,�w�1;�6ƺʫvJh��þ���jx^^D��4��?I�^=�4"�L������j�����MB���8^J��[���S!R�JM!"�E4"�T���	�/�@�H�6��	NĹ�3�m���}��A�Sx��f\}��������TS,����S�̃��C;@6ff\�n�m�:RG|�dy`\��2%�U�C���A�Ñi��&�gL��q�.̇0cXu�O��#1�19��]��Gf�5��Ϻ&T��'I��8��\��������G���M�J#���(�0� ���m���qM5�z���<�4c��MX�2�3��c���r��ڶnW�>?���K����͢?�h�Q�DC�� ���W5����"�O��/�dS׫�2A�8�+���i�p(�KWv��|Q��Z"�m%r>9nJi&�A��K���g�j�S!PW�@�x����}��~�0�1����a����`������`}zru�ي��?rOZ-k�m��r�1�B0;+U˸���ë�7��!�!�ߨ2�T�k�TB���<���Q��6��}��rY*���ཱུ;�2�nc�8�~:��!�����k@f�tm�2Lv�[&�16q����k����ҏ��
�. s���9�0�/�U	��ٿI����.АHYޒn���
���}�L�Q��`�~��A�����ą�G-�׊�%a�(e�wQ�l�ɥ��1 �-�E@-erKA�(��M�Kj� �N��>Ⱦ�uA(~:��?�<(*q�zN0�b�:�N�5��v^�3ՅY�D��G�2��ģ�P�D�#�Po��gV��ڟ2��{�&�!��
�������E��%�B���c���z�Z���j�F���l�P�W��I�:\&�	���z��}"c0[��X��.��Q�5�W�L��)<�m������Ľ��(q��F��N��a��V{��SL���(�>�T{�P��Z|#$6�/ke3�}�"[�3O�0�ӹ6н�"���R�pWQ�1���]@�&`�����V�u�wh�Ղ�1YG���D��RPƖ�:�p��b�242���I��|VĜ�I�|_�L�����	�6\��̱�3��X���ӂ�,w�x��|��P��}�NV��o�o� ���1�:
�K�b1��9W��K] ��W����ҕ���W�_�Y�O��r�Ve�@�Օ�V:���]&�X�mR<����y(�Y�w���1׼1>W��<Z���k�QO2�mU���.�0���{����ªp�Qt�mW3�#�^#N���A�Է��ޝBz���VT�*�� �X�3�~��8=LI}��zf(��RV��� 3P�.�BV.�/qPxɪ[�j�E�%M�Z8�r�T��}!_%�}���踞�:X1β�e#j��9�"~�iޫj̟��k��b1Ik��Ao�$�#A���ݔȺ�u����KW��eA@���cq��cTu�IZ�k�5��&bE�B;?X�P:����D���������%�����9���\:��J�;�--�
�S��hJ�����U��6��/���OMRR�����,_����T<�Ww��=+iyv6�ތ�8!���9����b�!,�}ʁ�x���L��怐��Gx6�^��a���E�["�E�r�{+c�Ug������=�a*��9��=l/�?�Y��_��+k=�C���-�c�����������!���:��#�J+�����1"�V�>O��:�T}xe�:��]�2М��F�u�i�?mӭ�F�Hs�% �_0����?g��;,q6�ųB�̞�1�|xc e.i�R Pu1��Ԣ����~i
%ܔ�}g<�h@�t���e�1��wL���F���0e�������~;ֱ��mP<7��?����	�U��� �:p�l��%D2���[�E�E*=Rm`��G�ED����T#�~dI��
@p+C�m�o"�J���+��ߴR(ͧ"2 �Y�<�� ��r�(���.�l�w
�1�9�,�"a�#	��eF��h#,ip,j\�iB�pF~bY������>��-j�:�8F3Q3��d�2E+0���WS��h��M�\�Sni�+�x����:�F��f`i!�ҸRVE��l2o�^�_}���wṺ�5�F���$$�&d�:�EHc�JK��M��o�����ډ6ң��(
e噮[�Ycp(qT�u����J'�>�D�����j\.sWr�|���zڱa����8	��sp�O[SZ��fP���t�E���QЁsI)+�����?/�2j�$F��жgW����MEr�{}��5ɕ�S�{C~;`��ٜ��^���R��F�	Ptz��b+��	�Az��:�
B��j��vf�/����M�����B�y��u���E�RO1�hj[>�p�<���)��%���9�GhlSS���U���a~�Ŧb�u}��Rz*{�jbW؂��_d��	����*���y�D�2�ׄx)v���ϙ�³5tX���h*�^B��O;��Q��v6q���C��WVs��z�FzEA���Z]��6#���k����� �0&w��R��yV�*�;*�ij��˥Q�"���|�؍ǮI$�]���{/�A׉�k��8�IZ�`��˓�7��'Ĳ��ǝ��`�����	�X;ў����º���d�E$
2Aѱ�ֵL=ɂ��6�n���j��a�S�����yeޜ�r�O�_FI���1�r���&�]�D�p�h�0\.'���
��M�J��4'tV��8"�UH[*Q���*�PKڱ�{{�@��/�hу:G�r!�q0��\5��!�n��R�a���氁L�5|�������ވNvL[j�V�q��먋���%^�E>$
b�g���U�oi�2�'G���B��� �L���O��s4/<��Z}�c��z2�<�Q���D�֕S4��2�gtMJ�&oܝ���b`��m�3��<b�J�]ƨhg~�c��zA��K�;u��lŘ�u���>�v���Tmw�i�?,i��W��tϴ� ���헚k�z(u|4.#��G(丑V��f|��T���M�#��kb��k�|/Cֱ�(�]�?��f1қ���|-@@�߆'�u;��4ҩ��d��� p��*��k��]7^�%leh��q�ޙf���
�l��ӤW����RwKg�%p��%�6�"X�iT,�vT{hMō����V#�C�w@����-�/k=r�V�Q�gӏ�.�{���~m�[w��W�y���M�{޽�姞Hj�W'��À�Q��̣Y_q�7&m�8�������5���f%�L��`����_RX*L���L��Sab8#��Dq���W!m��:�ד�6sM4GP�,�LVy�)�������W�]��b��X�2D�n~�
$��+Z̟N��[��@ø�԰��ָ�Ȼc>�fcў��hT���B(�\n7�s:��_&��7��z�Z��U�Sx���,�Z��َf_��OF���=�Z���;<�t�yi� ^O��h��˫7O&º��}=I�<|ql��]T��W�vJm����y[�w���p�7��q�*Su!�5	�DV����'J���mN{ѽ�R-��jx����s&SOL����^bYv�L%���Y��;�N����e�y�<��� ��8cQ���q�P.k����Y�=ݿP0i�E�XÆ�����÷�m���	f�*�NO����p+[�����f��MԳ�#��p�y?ˤKT����ܱ��L������e�)�<>E��\��1*	ћ�[�E�5.�Yȃw��ë�����߾�y���+{�^��rQ Ϗ��JY}��-�s��L!��y���-�wJ������#��Z�R��tpa?9�XN��1!\jv��$���!��^���Ȋ�d��DKx>�%��6d�Κ����9��Ԭ<ὒ�i�.�`��oV�LްZ�+����}�P��>ˈ������1I׋.�΢�l��T�ݱFF���פ�W���,���YXB<<�4�J�/&� �e+��?���A��.�Y]��z��v�G����3��º�"G�� ��*���Z���pH�� 9C���v���o"z�q,Y1� 5����BE����OCYϗ8ќ����I��S֩k�Cv����.�ZPk�/"s���kS��y��
MD� >XP4���\<���a��
O1)���.	�7R2��f��^\�l�DB����t^�Z�r��
�I1�wm��Rh|]�
 	�S��h�F5W�'�pv%�Ģ͸���B{SEk.\�E�O�̓p��o�܋w �ɻ�I3�ѿf�Bo?%���-���$�eG��z+�j%�C �}R�KۇR�7Ku�,��GC׸���=���������n��ힾX
�C�|�Kv�,z|�V��L�h�ժ�Ӵ���4��]SIe(s�\� ӄv8��F=6g���Е��V�Ģ�el��\�.~�X�%��B:��^����w��)H���/���H3^l<x�Լt�C��o旗��sӅ���R_%Y���C�r�R� �#q���̧����؏�v>\�C�Y����ƴ�����6���o��Lv��F�bY[?�[�D?��c�s���ʍ=�*����fͯ�ּ��������p�)�F�a��
���t��T���"!`��a���}�.�v��&��L�&P�\��2��!-�2z�{��Y@@'���Dk�	�=?�_`Д~*m�X`��L�p��H΋:,����@k�g\�ު�y�b�I��d�OWY;E6;��|0o̬G�w�wyi)��#��4�����l�u7��|����4J�Z���R��B]c$H��S]y�Вf��fxʓ����,�c��="f�Pq<C:��
��Ǟ7�����(F�F[T 	����۠�'�l"kNO�T�e�"�+�!?),~sIe�[Ԙ-~�k��b!�h�|y�{���l~�24��9���xL~��4��I��"I@^�����9���c�']�v�'��!|,�kݷPG�=~��)����'�E�D��)6�<	���
�O3*��3�ǧY��Kc�E�aF�ңs�������|��щx�`�s'�#@��;}˳fO'�}��a!�W#R�c��k�t �\a�ۍj�Kǿ�G� w�&�oo��3H.@��Svc�f�?@��Wa(��6���TOv�G�Nڷ�p�LI�\��8�P�}��3�;+�H ��[�3�z��?��V�Ϭ����W�~��'�������ad��-h*���O�j u��u7~�.�`�X�`A�դX����b@�+'���c�Ǐ�&���Q�X�� ����ݦ�˥����*��ъ.�?�F�]z-�A�ơߦ2��au=����)'�F��h!�m�ْ
�	M�#�VzI�G����-�d��k�0k��n�nx�x���˄�(=���\;X�Cz�.������<׫�kEja�"Ux�蘝܏��Ox���~��T-��-�5�v����P��X⮙p�
޵�lo$ni|a����0j�I�/|��n��|�|e1;��㥨G�[��	�g�f�.g�aɑ45"��ڏ����B�Ʋ`��s9��.��αT��;Zs;��8�<}�(��*G��1�`�F`�� Bx=�;3�d�0��\�?՝��iϑu�bS����}I�!���H���@m5?���)t��*!���vt���؇�ǉ�F��<y�E�pyNa����RW$�;��?��E(Z%'a=��x�Ǝs�]WG;���my`����n/�:��Q��M�GP�����lS�l^?T {��L1��U����|EXEY���q��e��]x�[(-_���k[�p����DN�#*�<2�_����J䂁�~�L��ƚ{T�����䍙3:�U�
1�t�
vɞ�uJ�Cc<�n���?�l Rl�� ܺ��A`�����8�Iw��7�0��~
�/˂�ig�p�;�Eą�u��&��M��h�u�?�G����O/@�zYƔ�ϕ���]sS$���L[@���S��a��WǶK�v+dFH�I͢#��(������ֹn%X���d �W
�7u�7ߒ^����5>ר�^N� �YR�A�S���Ae6<OTI�:Т�k�b��P�?"�`�6�&�����5�����yL�y�nx*�M��4�ԣ
v��h7�Pg]�hck�����c�2�Z7�9�vn ,��	�w��1H���a��ZR�KOSe>AڜǔAK�K��ť�[��b˱��U��Hԁ�Ù~42�@��;� �Y���
��C1�'��+�x����>#H�b_)"g��wf�[�7��o��=%�����ea��gp�\b� �/ݷU�Y��-� r�sgv����|O��fx&���w�D�����8�=q�]q2,��6���Rr�]B�wY� ��r�	Uѓh��{��R{��}��}:��% ���*�SO�Sܵ�8J�"�w�����)˗;O���)�û�N��xK����V6yu���0��0�Y?����}�4�h:�
�{qT�w@V�iy>���`�Y�$r����Y�Z�ؕ�A���6��y4_h�x�M75u<���кn�p:�o�ke��r=Q�ȗ�~�*�'}�1���C�7��h]�2�md�_�T&'��F��f<�H�����[�(��L�=����B��U�d�E�9Q�0�'7��R�;�ˬ�Z0ML����S��><���K��l�m
�d((���)��/.̖N�U���Q|@�:5�9��h��U}�	�v���?�ꮶʟ~`�tĚ�B��kP��6������X���UlHH>���H�x���������HaJ��%0�����Nv���N�g�o��ՖH��,�~G���^T�ˈ ��Ν0�S;����BZ�����4o@c��2o]�\鞆/LN�5M�QF���|�A\;��`�j���*�H�l�X�k|�lWC��
Ot�r$�����`L�&F��f(;��}�_	���2�nx}�`�c�ξ�������5"]�e���&���f$7O��~�,BY��k\��3w8/�AL�k.<"�bY�~eu�,���G���F�����?4��i�'��`pY���`�{���(mF�.`h>U�s}4��#dn�ct�L����s!
��L\٬?�@�c[�Byg���T`״��M 7��$4��^�8΁��6�ޜ���YAS�41����o��{_��:��m#�3k*��F���G�^���_�<���~z�j�L�-D��e�qcp�͝M�s9���b�p�)�]ay����9��h!�:$$=��)r6z�zN��T�G��(��l��LE�����#��e����J(�ʣsXL�&�
n��а��"�v9QS�<2,.�I��dbM����0}�;����}�8�K��1���M�=�}�/L�9��U�s$���b !����jr1���f*w(�0_B�D��,o��\����I��9M��4�8���XLH���-�c2|�׀%��.l��ۨj�n���ԉ8�n�˲�5�h�E��^�آ���D��q��;NmE��ҳ/)ROǳ��1��.����Z-�Xj�l�w��iC9��������8��;[=�"��/�%�|M��}���aey�����^K�0�����WuNEX�f�
�j�����ֽ�.���ź-�v�\�����?� �Ѩ��vj�!9��k6�ɣC��8��Q��w5�!%�M2#�_e�jx� �<��k$%�Ф]�Gꍖ�j�t-O�;�^xNH�|dO��R�%}�J/Ý�0۩�g	<�%ҥ��܆Y�[FM\��X)6F�l��F-L�^��[�|S.&a����|<���4�JA��q������v��-�P�3zic� ��:�����B �v7��ğݴ��H�M�2����f�8,��2�?��%��t,y�c6�P�z��G�>�-1��W����
�o�n?����3!v|�-˨����׻�ϰ�;���oNT����u4��'ıH P��`�|�8��A�9B��}����7,S/7���7�G�!ͣY�slI�4y=<r�]��L�%h;�K�E�Y�o�e�U(��[!���.r ���Є���7v�B]LW��E�R��#�N-���rz��"��� e Mf��xu	4x�G,v��N,��J���
����"~'������NTn���n-2�1Nh�"���'�bO��..	*���]U�=d�
�y�G�NF������u��O�y���.Pz+2��"���+�i�%��~Jt(;rw�+w%���0M�{ML�jA��h�?���^�IEꎅ��N��X`&��Y{������'��b�*|A���!��/�D�%�sHG��&��9cD��uk{�	S�ϣe&*��U:y��o��G���}~��@pC-��_��F[�yՒ�'(5�i�..8��g��:A�/��_�"�me�>�1��`�٣�_�%3���S\;G�%c�F8��$�/��f�:n琣�-��V�u�8�H<���4?����2�~�y�����W��j�iQ']�Ɲx����?��zP|r���j�����NY�f̆�+(T��%��:J�a�K3��w�?����~�n��M���3]����Q?96@�+�B�b��.����O���d������kExX��Ip��y񱯛�#�J�~t���`��i��X�s�&�S*W�kP��n����߮Z��(���>�3����T>���_��o�cHEH�m���,8+j�����r\��)Ζd��m}Xc��&��V�MX0��"�K�Rp�!�����{��|��$���}Y�S�tI�Y��n:_�����p�R8��������mКs/�g�"��+���s<��QfSo����.�-��� u���Ԏ�FBn;#eip�,]��������,��E~�����7�?䝱����u��zZ�d����S�v�<l�Ͼ>�[�tP�#��=P��/�3El��0S�����T���_dɧ��$�W�7iV��z$�/_m��"�xd~�M9������'
T�����3c�F$6�z�`y	k��I��)����)�U:!��n���VO�I�$��,���~ �c+$���F,�Q=r�d�eY��R�I�G��Q�G�յ�.j�����}>�Z��qJV����O�$�s6��Q�`y�>���h�\EZm����c*U)�ƉB�%�v�Չ�z��̲�0YG�P?�����*X�,-}�=�m�@�PCƎ,?Nl���*�y�y��<s�^>t�v|��F����h�g�q2��_�M���A{�n�n����!Q��X<ԅ�=���[%����0�E^?�~�@�_��[��eRZ�]���Lc��70���)�؃���>��a[����.˗�_�qB�+���VHx�u���/�Bi�����2����A�j���Ǵ����]��I�h���d�|�|�������OGQ*���mT��]�-�����x.8�U��3��{B���{Y"�����v[-��Q�|V!�S@{�s�c����d��l^
G�bXl<�����].��ꬄM����Ԥ�t���g�Ĵ@E����{�Wƿ�+���?����NN��]�3^������G��CؤK`���iߛ���ȋ~2�Z֬�T)X���s]���+0"���06�G$N�}�
l�ݫe'���|����a��D�\����mfzIh	���rwWb�5�_�*�H�c~K'���+�r�I�}a�T8�K����!0~;7�8ʦ{�2���i����N$h6���;���>��)~����%]����c�m�}j �'v$D��Ї���|ј�e�
��Q(�ßF��{��&�m�}	i�z�(��UV���%�0\ǰ�wN�`��:�>� n�þ�Xڨ�
y��PiW���)l}�LDE� �&o��B��)�Q%OUج.@�7ϯ�s�$*_��24�pԯPԢX�0ˆ����N�V�!�����|�h�ݍ�R�H̯Q=!�O^ؖ�)^�����T~�߉���K説��*�Q���Iw�E42���� z�V�0a8����Z�ǵ��4ܬ�� ƌ飾�b-�c��@Tʪ1�=oL�kW���1T`v�-�+ ����LрZ�V�dAB=����\�y�ȑ�^[_o}�,(f��!��U���?�B���Ã�<���9bt�����d�G�l��υ�y`ՔQ�O�a��.N�YoTw�u��+��(�3`�˻f���%��[����5�
��6b�7(02M���4f-MF�|�ޖ�cW��n�8ӌ��,�1�?��bdxJ#?��ץ��SK�SuM�����
������Nn4}C��Jx�q��5Ftg5a^�:N7σju%���!�䠗��N?EC�n1ݜ��_cЧbI�1� ��a��������K$��;��$,�"���t'�b2�����!UڱŻ�m0LA���y?r!��u�$z�$�;���W�5��r���Cz�e�ऴ �\l=d�c_Y�7/wOx�������e���Xl3�S�m�[*"����L�y��F6	[���>��4F[�O�:'��7y�1�mh���^���9������D-ji� s�1�hg"��!�,�6���Y�d�c���_b�Ȍ%�@�j!B�KD�X>�o7 kR���=0���<�)3l�k���'c4a@��ߔF%���P�6�`�A-pD�>."���e���D��vi�C��N=kb��#�pǁjt��4޽z�sj5��p���O'��Eҕ��L"�X5�r����X�4�91�;˺�͉��n����k�[�kSE�{qr逐��B3�J�����M%v��a��{KBPN�M�H."�KA*>�m]m�"�����.��PJ�K�!��*�=Kڋ@s2%kr���o�$�w���d�K-�_��2Z-s�ҁ�.+ 6]�M�̥��j��K�L�COX~Ю�b�Ԟ��>2Ӳ�.�̺��A����Je�as��oj�&�y����u�������	/ˤ�	� ��:���ʖ"����"�3+����|{a+����fm{�����][��ptoe�޴��7^x�eD���ƀ�	oXnf���s���x,�7s����py+y��o"��iw���>�<w���K��9
��\�@+����_����p2w5���;!7a��t���f��xP����<@? ��*>�Y+���2mU�w�[}���hƞ��< ��R�Lf�q���V��N��2q<KF�+��η|�_����|9�|@l܈�7_*��eU�2߾���&�;���q/�C!�gI�V����{F	��r!���Fy��\Qb�$�)���_}_ִ~-8��4��G�	|�`�柯���0l�&�ʽB*�QE3=�曛v�X�%��_�Q����%��X�RU0��[YyJg5aN���� ��	���4f�����;BЉUng/�F���ШM��&N�il�����q��O^�?e��n�k ^s�V���	u�4�m��f��uϕf������^�v�Cb8N� �4��p��19�a3_9*���Y$y��䲠�$6
o���29��i�Mq`Dk	�L��j)��z�R���l��e�Է&�����nI��S� +X� }��̞fD͆�[A6YWoQ���(�z�����j�v)]�;WE`��Gb�K��&�K,G+jYN��,�3�L+���gs���]ͱz�USI.���ڰ������4�S�|����r��!�����A�d �&��6�=&i-JuD������}h����D��	G?	�>���z�2ni
��g_�U�@jZz(\ͮ7l!3���=�M���-�tM�"�b�}ܸ��<��]�.^�b�]�|*�Ka�M�3D��)w��q?Y+'�L^Y	�ƨ�g:PR��Ͳ�/PN떴�F����=6���&ɦ��xB,��������Ƃ��
���)� U��w��������Xꕅ=�<ޒdc��aތ��RHu�9k���ؖi��;�g͇���Q�?�W�]�kbv^K�ݒI.����%A���xYO�/��P���V���aIB[Àf�[�Vv�9YT~�F9�á�liv@�[MA5՟��ӽ�EM�Z��AKg�;DAZ�cQ��Q��Z��d�Y�KZ��O�!����y���z#��G� �L4�S�����M� �ӆ5���QA��[�D�n�)�o��?C��lѧ֙��bpb�S���6�%�u���[�Ԁ񦇴pz�d��������ǽI�d�[��ˆ�7@a<�����iV�ÛHZj������b��,�-�g��a������|��0"c�����t��/l�	�\!���'h6���b��1�N�jD�4��P�=ѣ"1m���	�h�%b�Z�\��-��(x���%����i1�C1?,�P�]&)Ds�Fc��Ty��Y(z�ɺ�R�ٌ���}���,_Ũg�J!�ň��,k	��?��m�_.jE��׎�F���OX�o�<�?l��Q�O^|̩�㑝���Z�p�ϧ4V/����	��^H������L�<�+:B����o��l�rg���!ͨ;��Ҍ:	�����/���2J&�hO=TF�W���D�3��-}!;���%V@lG���z�2\F�|��d���e�G�w0��vD����0�m�����2��˶3�Ŵ�U�&6���H��s��)�(��xi|�7ʎ���$2H%�����2Tw%j/ڔ꾿~
<$8����\0���@��u�&(�\��_on�E���Qt���$��[|X�����A��7
:�MV��*�}����&�8��EN�ī��G>5w������~��� ����E��74��h�L|�~2��eG-<~�C�iB�5$Yal�k��f fUmY���+E��2�����jq� D��/$�.pҤ�e��+�I
/*}�/��6��Es�
�Tb���[�fYhv��|���1�4p���� O:�f�� ���y_��iӼ�p�J���v]�6�w��n����3N�K��^!���(��v�;(��d��ʺ��E.s(�o��Z!(%��vh_?����锺E��&È_V���q�fh^�
:.FQ����Uۯܜ��>�2����K��ôA*M/�97_���x=}0�7�7���_h4R��J�z��\�m>^�WB{�P
�{S�p7z�����I����@Ac���z���ޮgT܏Jh3Au���3��|G��k��ݚ�X@!:�+���(����xZ��P�}�s�)��/I��W7�-5���NPfi���^	�ϷE[���5�BM�y��1�4 �����}���3O/>bR��8�x�(U)��6�pv1`x���l)&>9�%� ۹�q�4�*m�es�B����y�g�����s�[�Xd��	.��ϩhͣ�og�B+B�Ƣ�5��#������}M��!>:28(����_�%���B��!��7d�Q��u�I�5�$��J$x���}s+t'j����Gc`�'���A�������/4���4>�6���8մF�gX��]:�ȯ5�W����s�)��瘅���*�R����N��P��oZ��7�4��W���!�eUmE{^j�U\�t}��KTD�;�
�k�O�)����/�� n��@�Gy�,��L_���P�)ǆ� �4P7�|�?EkE�A�Oa��R�}0w�7�CM��7Jo��!�C�����a�nP�H�.�M�=��q0�$9x{�e=�i��.*��i�:�C�����9�SE��H�̟(�.X�� �r";N�WW2�7s�i\����wt�1Ғ*� �+dNN�)��(�#\�`r�vv1	v�e���2  ��͖����P%yk3���$ˋl��ޟ����?vz�vc�W�،/��'v�>+j��G����u=��}��Go��P,��M[>��z$z!2z���m�XHo���A�D� ��'@��@ʘ���9Q]�%:c�5��V���m�ꧫ�$��\����]����֖X������t5K0��Q�,_ ��n��q�}5�AF����q3��C=n4�N+�	�_�����K�s�ӡX��ҝDU�� �ݫ�B��ÛNz��������4~1��¾�N����a7T_��E�-I{�cI2�V]�E^H��Pt��!HcJ��k��Y����7�t֢�~$��?������@�c��oHx���צ���%G^��Tqz�׬5�>UN����@�W��1pr��<P�P��g���MԽ~���\<L�b�������H<@���Hi+�A�u��ˈ8��ʚ�F��U:I�����z��C?�[����ZWG���J�T@�K���j/�A�גi�i�i3��3�3���f��`wj�Ӂq��HY�LXk�������#�G�U���0����S0��WP+�eAR ��H��ا��� �������2�2�I$�����:LO�3�o�۝7���x�U ��0�6[�L�����HZ�f�+9`DaS_�I+�\���'��*)]Bj\�ỷ���r���\�+'�^�Lf��(��0m�_�O�F�'V
�Ss˒@��os�I< 1ի^'P�����	� ��&����{2�� =|k6m��
Ǩ��IL �\�qiVX���S-���i-�c��a޿�Q��x�B���$�T1��R��M�F,�{+UA��v��#�	jT�{�e��/��]Wt�6���t����KκBd!Ux��#�Z�Jk�#�y�Ҕ�,cV,�#ϰ�8u�9Ĵv7�0����7bs!���R���vb���Ǵd����[�i�m�+D���d8��y<sR�����[�0��8{x���oq\?�����8`�]����d�dL��ɤ�F�oQE�2 <�.�^��6��������=�o��d�������w�k��w-�Sp�C͝D43�`�/ਸ਼m(��2�Nŀ��W�J	k4�)M<&�$.|�?�����"�$p���Y�].b��3a���>$��-��8 {J>	|.zW��7-�_Z�(�������ˇƠ)�D!>�Ȥ�
���#�w�ga����b?G��%砡}�N��Nc�3�T�yd%���?��ڎ-s�/�#:9z�}�5��\p7%!�x].h5��iҟz���EUl�
m������~����U..�]�z��yS&�,?�?-��I'o|��|�.�Z�V��	�F]L�̂h��-��6����>���41��K�Ѩ���/S/F��*��̛ ��%;��<�Z�[��!^qH��e����i��t���Y��r�RCH��Z����	�r�/���5�/�L�D����y���"��1E���o�V�}����n������+Z")�}��/A��{�/�y�t��%����=�8!<X�մ!@,���E�H��zp�9P~~����
���Ǧ,�����?<>J��5/r�w�Y^��C�r�5�X�U�;x�\�9&ϿCz+�0X����˺�ڬ<�x�=�~�-�gB��k��U�<!wU�:g��ȏĬ�����qߏ?��|��}�4�Z��T�Κ�='0֙O`��'.�K�ׄ~ w�6Rv5�Uy������%��|�
��X/E=�Jmw!��j�0�?�,^I��6�s�Ō�]~ѴMЙuč㑉g�F��mn��U�KS������F�m(���%���_�#e1�z_c�`�Ɗ�pa�nW�4j=���G>�������W���8�)a��L��A')�-���&u�i�z�!Ȥ� ��%���F���6~XcB�{��N��;�O�o@>���Že��Fӫ����pyNQ��ɏ�ߴr���.�E��{j��Q���6�2F��e���!��
Yx���W�_82�j#�m�y�>/����PSS����t���\001� �7�x��}�%����O@�zrt�h����{.�A1�**c����#<_V��ӝ#6��y�J6�28�u����~�I�ϯ�s���yERgǎb��Y�C����J��uy6����b�	U}�s�}��*
�1�g_G���B���
]�,I�u݇����W�1LE�oe�W��.<���N@�$J��X�ö�|�&�V��{nk�W� +T���3�����A��͹`؇/+6WSM�?\��n�=E��.��pr
l�=D?�p(���y�������rFU�i	p����M�ބ*e"K6D� }5���j�'_E�{!���U����w�V%a±�:(�U4�W�i���|���㒓��hWH3�����%�ݮ�/Nm>�����L��
��W�����%b�{ֺ7K�u4N��{5����"K�p �M�
*L�m�KQ����S�.��_}-��ҟs~8�x%�5~��`{5�уY�rɰ���9`��)d�N�>��zp1��x��H����c~�q��4�*���6�Ӎq#� �&����`��h����!F9~�����?� Rd��e赿+p`�W�1�+�}�^�ފ��l�k%��_4D�?�T-^�7�`+{[E���.�ű�{���꾈:��F�9�k�3�a�faI=��d" ޭZ��[L�B%Vp �x��?H(�C��)-������\N'�w��;���"x!�ը��-)\w_ήΝ(�N�2i���ZnH�b��v����5T���yW%R�`�e��Oe����s���yH7"����\��@��pŠ+����(Cx���+��|-�}5�8���վ\�ΧY�ˎ&}���b�1݁���Yy�\o��_�<��ܴ����4M��D�v6�%^�r�Lbo�g��l�)���>-B���  6��?����0@�@̥%�E�*�����}�]����4�&F����4}#d!ϳ H��G�¦�J�SV��PG�#������{��~�<7=�X3o�n$���C ��uSrIag;�T���r%� ٔ����{y�+��H6/o2%/d�wT���3< ���u���xy��7�K8����շ�J�����9 y���B�i"�U�����p���Lv�h0�xH���-K 4�Vs9 L[4n����.�OG�Ε/�y?f����X�J�[oR�E߃Q�����NI!���K���h|��V��ac��� �s�Ik�\��>?������B��_����u6�&�8͢���kSHX���yǲ��I�!�S�[^����0�}�Y��NfԖdw�l��)r��8��\�����vX�}��^��2���TڿiZ��]�d�/Tk�����n]�ש'bYj��t�(��%����Ho��z�P��B=��vZ�}_+��E�Y}�>K�n0���O;�#Y5N�R����h�l3���4 	�2`�z�dGֲ��ͭ�?����\(�����ĩ��@Q�&�x6�k��:`#���{����f���ثb�Q����'�f�I��5��N�nK-8u`1}�m�a/���������Gpq+4zs�K��%���HD^sS���o5t�cA�tE�VR��7G�N�3�J��ׇPOV��Ǫ;�9�x��^�g}h2��s��u��y�����0v�m0��Y:?U�����(w��f��:�b��C�_�ߓ�zI�l�BfW8&��ݙ�*c��d��Rnw����`-F�� =��x��^6ҧ�$�"���^>�$�_O��3��=1d���s���W~9�^q �)i��0�/��W�!��d�q��o�B���IN��J�<�cԬ��Y���P��q\�B�]Ih�v�0�7��t0+��&�Ww��l䫏 ��������ްs|����E���U�2����H��Fv�, d��0'>�!����Sl:�Ŝ��{�v�N�Ѳ0�G��<o*-��uFp<�����S*f*�(tᠪC�<��[�N$�l�.�z_�f[�hK�>L5��[+����\k,���}�=����ͷ�L�\g.BM6���r�>��NixG0�����60�m�jj���T��a��qt�'G���U��7�]_�(�+���G���*�+3 v��X���3�X�~���o��p�$`ri{>0)��ه��J�(�D2.��&�t�g�L>�kf#��n-yhc�����_p""5i%�۟�1��݆����՚d.Rv�I�eݖ�}�������>�t����T$ǀ���Z�&��j��}��������>[�lB��hw]͖��]*�+%�B��OV}=����]�|�;W\�J^�hoiQ�|�41\�3��(��S��V���@�i}���7fz�ݓӟPP�0��!g\	{a�����o��1��m�	<����O�p��w<�#��z'�Y�{`�x3�@�%������ⷩ$~��:�%`KP�dE�?z�� D^@3h��5Q�'J�aِ�=�o�$�X���KX��YlrZSۊd�=��P9e�%�I�����.ǜŅuC���p�%	�,m�D7�v��A�Mp��J�ѻ�y� ߓ��m�	Q�����z4�&	��i?p���1fs�לA.1%��t�V5�X��3�c�����l��ϸ�-��:�/���6$�$��ǥ�����p��Y�N���5�LԜ�O>�As��b�!��{c�%'@q���Ɍ�z]��("up�gBW���m��U�I*�8�蘙 �)���a�p3G
��P=�Oi�m.�����:}Sy3��Z敀�'LަDȭa�V�Zs�+j��}=�i{ɻjUG���&ո��m����e�&��)��4��y�
9�m?,t�!�<���ج�d���^a+�ɛ2~A���3��UK17q�b2�Hz$���:/A�+��\񊄟}t`V�^W��%��#Y�1����qY�?����A�^�Wf$.�:�Ƀ���b-�h8Q��A./�z:7w�	�u#aH�.�P^��.�̸k݃����W�������'%*y�@e�{״f�}��y^PԈ��,��4{��$�F}��՘���J�0��R�uM���Kʝ�HNz�L��/���G�,<�r뗿E������9a5��"hl���d�iO��>bt��)/η?/"xٹE`�>��t�TOB%h����f��SYn`eg��ta�
�)��v��v�XC,>��u ��S�*I��ubG�fo���n��Q�֥����x�C{����M�=B�(�?�:�S��L(������rۍ�@f��;r:��M��I���*�����P��\~w}�z�	��0R܇,�q$�=f�XU���tk�=>���e�0X��,tj�E6j;���|<h����#�����-�����/_���t�YQ����1�yEP�2�M{�3%�v�/��6�:��7��������o$Z��"��������c���"�tm(���u�8�hV�����;
cLY`Rqs!͂�KL,�N|^�T"��y���i�͒��h�ߺ?��=�{%�o�;������8Lz���z/ʑL-p0���A��P�%����v,G!��;g��˭��T��:�OE��s���F۰��M��l(v�1�D��o�L�q�7�i`o�Ɨ��]7^��z�K�φ�l5������0�l��c�F���y��k��� �kӂ,Eb�WCc'���`�Ȃ\oW��9ޤhp@��K�^�yrq����4RD�?g�-�o��Ȳ�u���!j�nIV�Nz�`?m >)=Tx���u9�6U�֐o�w���1������i�5�x'*�Ok!�}^������X���Y=S�د�Ʃ?��ۙc��DÌ�!j�6�@��'V��R��=��j,�5�[@�!v{�;�
~����Y�¾�y�A����u#�k���:0��ړ���u5�L���;^s:�^����V�.�=��"K�o��OF*�T��keD��Ф\�"�����+��~��lC�Yx7ϑ��c5����hJ�]�%]��Tʱ��(�L��Tc�c��>�F�(U�>�
Ӑ��4=�%u��{`Ig;��o���$�T�Y8�p��X$ ��
�x�j �o�vӃ3AiJg���l�M�J/	�� �g���*ډ6�Rk���e,�RM�n�W���ƑD�D�fy� U�ꏘ����#�<}Һ�@{��Ә�m��mc]}����Y�t�Mׁ����	.=�[Ag��@�	�3�r3
�8]��Ib2�f�2P�F�W	8�,w�/KHR���-�1ĝҿ�P��l�'��!(�hQ��`�g�zz�Jꢪ�1xI�A���.�3+hk����d5����AP+5�G���V�^L��h����R��X/�E��^�l�yS�e�r%� �p��'���&w�޾hɢ���-;��OJ���d*�t�F������9>�Xɔ3^����`O`]H#�9H��2���E��d���L_D�w�B��ǫb-��Z)�����u�Out��\�� aY�l�`/t���a_��h+߹��>��RvV�~� �q	~�W�S���X���Z��8�/�2D����Z���,�dP���2ս��<`�VU(E:�3��#�Q }�0)�̳�np��a� ���{b��\T��l¦�
@�Z��g����k�]c�tv�ѣQ�����o��+�F4�vG����0�$H����	�]˵��c�U�U�1��ܗ�J��'�
_`�ڭ��`�� ��A��O���}<	jjN(��Du�r�`�%lކq�ߕ����2ך:PPq�����7�.�I�8ii��J���/'S�88<��y1�M����<����I��=o�Z���
P�0\�ġ���(�Zc@�D�JJ�tB�쿛I���>���U/���tu���H�#�N��1[,� V��s�N��v�C����;��D)���,XNj��&�2v:0�fX�0���_��L����Io �`H�l��e�F�38Drӂ7�҂�����jA
�z<U��������Ԃ����+I5*m,D�
�2��:�Bzn���.�WHJ?�׺ˋ�����g����i�#�N��Vߩ�?jM�<�4v�"D2h������_\m�#7�A¯��p(�}@zt��:��nh=�*n�H�3��n'��V����et˥2Z��.,D �����);�`Xz��qIt|. *��*����o��We<��"�ػp�����<vV��(��$���|�g����+�'W��E;f1��z��K�����ܪ�Ɵ��
��0����M}�1Q��}Bc�׾B�B`g����
��v-Z����(���_��j(4�L��m����#�ۓ8�*����!xպl'��x��/ƚ ��]�ǜF��{)Y;���h��bdW�~X=j3{Td��* ���"�i"o�z�IniRP�c�
�TE�L#1@���*�u
%��?`�^Nrz�!7y�O�����9���nX9���~L[�hN2�@>�j��q0��0�ce��A�����3H�:d�l6�gG�2G��I��E���f�]vE/;���&T������O�� c1�h�)�"'�=4��ćt�<F��帀�dB�3�C�=����a�&z]g�ʟ�TҒc^�V�zX������a4��YkW��J�w4��h�s)��v�G<�ao�t�����Փ�/��e �к�I�{���7�JptR2��ZK%�v�������;����w{�B��q�|�l0'J�ϗC�e>5�Qw���`w�=˫QmI%���}�,_ޡ��%s���Epl q-�_���5�0|���gND���+mKU �\��oR��"��i���qZ����L-U��_d�Ԑ�^8��~&�lz������Ъ���-"��ե���ީ�����(�Xu���V�Y��o��Qz���)R������ꔍ�	�����x�sJH���4k�^4��^>&6$�9����̕�an@2�x���K��d����;�ޢ�bzk�?Ŷ-Vp�]�j��`�]�hB�X���)���*5��).Ί�&+z�*��uݳ�+5���
�l}b��c�V��6
�7S��Y�>&�3H�X�!�P>6z���6���,��<��,93"���2�g}c\��%>vv*P7�x�F��������1�>β������2/�'����͐0�tg��b_d�õ(�)����J�6��V4%�l����zӌ�T��ca��Sq�y��_����	{�c���q6%�k$�h�x��l~�Ji�p;��o��0D���u�Q�ߝW$�B�N$��5a>Q5� ��;0�%Rk�I4�����ɩ�'%<y�ۮ���朡{�kK�}�^C�4Q��ε�<iw�L�4�Q�^ae=*_ku�,s��]��L��1F�&6��2[�"O��*�t����S�k$�P��#��Q�
���-,�����U�Li��n��+��8�SGGE������5��}��K-b�_F����9&���A�r��aȪ��U�d��V����M�z���`�	�� ����B�NӪ*�}�D�./(�&]0�6��`\>i�׭O�/�E��@w�2f5�8lO<�:����`���B�+����/�ic�ĉ�5&��]�����;���	����Xz}�e��ਫ���}K�x\���6�&s��9�;a�|)e�,�'�C_�y
�s�Ja�9�
����'�R�� �jR5=���8pGv�8}cg�wx¢C�!�SrƦ����M7���<�r��U\>[N���Nw�u�/-�/<O��-� HI���$�"� i����	�=g�J�A͢:!��Qo��A���^����� N��Rc���<;�_޺��z��^\8��L�.����Ph��/zm���b�� z,rI%�I�@��
aP���%=����y^a��N�z	0�P[��S�
��~�|4�5[l�tz�!��Y1�|��ϝ�5vkƾ�q��5�[�-?ﭽ�f�>���&Ձ��?���C����<'�/�^� �>3Ӏ�?ȶ�!�;���N��XG�!�
*��[6�r�+z��,���ӽ�l~�К���U���"7~�ʖ_���� L��S0��I��)��X�Q�?,r_u��Ӭ���|%ҫ�/c����yc2Ҁh�C�}�Jq�]��}蘽�~���3罿}(}
��/3��d�9� �ˑ*�D?u���<�C�x���}.&�1���rߪ)���[&1���PN�B��҇��L��U�K�OuR<;sI���
Ձ �l���}՞&gU���m�,k��I�vfk�����C�F�+\������s+��R_ĚlV���k�?�a�������>����F���K�/!}<���*H�x����S^ȳד���g���Ĥr�ÆB{�W8/J���%�C��2n/Ԟ�|��jb�6��ڽq�DS�ND7��=��R�Fԣ���)���ri/�/l,n��hn�z�1�s&
����_�B���m�9�ΌG���}��S��>݈�f���d7Uy��z���$�&H��Ʒ$ܢj{�pW.�Ֆ�lJ:fS�H�j����Z-�!��ȴ�*�t��h�Z��F�=����,���M���~�5��9
��,��w58<���s��/��i��_;�U=L7�ȅ����P�'{�".�yi��ڇLG��c\ė$)��G}��/D�a�tGo��B�a��i�~�s��D�|��q!V��Y0.W&���Dht�^K=����-2��A���hS���CN>H��D񭂧N؏�*����[�@��7k�?���)(��v@�����F�oR���OLH����%F�4ݹ㛏���et�0�*)�]͖W~|I�Y'�@��ГI��$T����t{P���8&��c�ͽ���B&�=�4���!.�[�\�3#ܝ�s(�����x�zg�o���|��8��>��H��*x�����ǩyԈ�4�SF�J�")�?�bn���ur����m������I��e��/ή�>�Lm��Oˆ*�1b��0YT�����V}o1d<v=�l�0��Q3h���f���7�`�3��$L3��D�0��\�7l�ca>\�wIv�I����n}��0b.{�(�,�F������9�W��A��06��[,��6�4(�B}�r��9J	�\mI"�imp#A�t�ݰ�4w>wσ� !��F������f�ⷺ��p���k�?�ԫ�dE2�E��)���]�J��,B��|b��Pm�"ϗ��$-�#�E���e����d[�k���Ko�=�܀I�f�rk�p�oo%p��\��8�
�f6jf��X�i~Ma
�bGɔT������aV�)��"b#��Q�4�I@�����^� �Q2PTĉT�xp!�-��=���c��;6>����F��j��U��ô��ӳ���l♕em�.Xv�}��j��0C��wa^�ߡ���*h� >0�q�
�2��ĎUp���A�I�J㩊����Ӟ�a��R�a�W��"�/v��㶮��!kSi�vqB_-�,��� �q5Ӝ��H�)z.I�Nh]�t�i�@/����/EQzٛ��ō��L��e��I$�b�)�3Me�>�Q�0$ F��	&�4�'?3�g����,ޠ������^<�2c���Q$����m���jyزW�5��!U�Vb���R~L?��̒/k��n`H��{'��C�ؤ,�w�ԟr��#-$�����k7Z�3;N4����uiU<�L�=�0R;�jv�*p��s�DD�s��)@3Ϻ��QN<y�#���[�*���c����?M�L:/H��T��ǎ֞V�ޢ�C>Q�!)S�ȅ��z�"�;qv��[2\B�c�W�B*/�$�8"w�DG@�*Y�� �LQX��)�]�\Sw��N̭QXA̓�r�E�ƫ�F���ES�/��s�[.�yT[~]��-�t�c�@�������Nm�J\W)��Yp]�i�~),���*.��A��ێ�kO鄥e��'?Zt4R�,x�{��#�e���n a2}-\���Tګ�R����!�k�#r�E�W������~��o�d�QS���XgP2�o.�=���y�΃���j�C��C�v�^����l�Q f̦k1֚�1��5a����C�)���v�?�;4�>� :�tQ@�H-hj�0��z���4����::���hm���SX�b�Z策ZUsWv��L���wXVl��ä{Ux��������_��|4���R��;��9���Y�\n�1�"-�����%��a �}w��\��敂s#�.H?'\��y!�#BO�l����?+� ��9:y�Ϻ��7���A����x�V3�O�v�,��]��>)�1����#�Β,T�9;�	�g�b� �'a�C�yLw+D��r���d�F)Y�0�A�����<�M�T��� ��C�+N�B~�8�	B3�(����n�P��&�8���9���0��0�L@S@��2Ä����3P�m��_z4J�.f����2�*ű��p��aa�5���s��P��0�Ϗb�2�\1��1��m�שI�2
s����xBU8قpD&�d�<}6Y�&�w4Q:�w�)��_��f٭�
�Me�Qj�^�']2�q���Ә��x���~��̈́�E>�io���rODThK2eM��yz�>z�Vf��A4�/�wf黝�B�.�|4����Mn���vp�\tL���V�e^��|�beձ��մ��� BbL<�����k�$3X$�b������|���'P:S{��M�l&�f�$�2��I�b���G
=�Y�^��j���T��d,�χ��Z,�W�9�{�����Z-���B�9���_��s�ު.���%���Ǧ'�5I��%��{���;�Jzߓ�U�c�^c���|��� ��d ��TJ�5T�e�@8�%��k��(�t%�=��1���;
����-öb%�MC=]�H�8��}�F��&�#Al�]X;�e���<��a�j�U�=���J��EaLhN]&K��߿pQ++|�.loGM��>*!�L	�Y>���5�����$�o�q��T��J��U5
�z�n�5�~�%��ms�on���:�,��M�B��k	�8;���MPp#\BgE������N��s�.���u�t�"�"�iח/ ��v9er,z6��A�/ׁE��O�7 ����ĳ����2idL�~1�ڟ�ESf���5�(�����`�]���1ٻ:���X��%�(���{L�G����?z ���-=�4��g�B��%E�E�[�'�ɨN~�Zy��"]߇���!1d&��ԁ��`�F�v[���&YY�߬�3�~�Ȋ�v�NW����R��2�y{!k^��90�7X�sTe�\gL��_%�w���,�qI��c-������?5K�F�ŕ.=c#L[�.��~ޮ��K�Qyn��n�Vq�K�|�:�	d�JC*A����[��ؙ>�eVwY�i��E��U"��J1^�������*ܿ!Q\�������Vd�ǂsC����#S��؝�ބФ��3������@]�Y?V���jZ���������q���5�c�@�tMZ딽��S��>:C��]�^%��@ʑ����~�����Bv����K#W�x]]��5���
WɑM�5,$~�=�1���Âw�y��X.@�T�ah��M�2B��̖QH<X�辈$o7o��^8l�J`L43��y:��p�������ˁ�cJq��~ff��n�g�R�P�(�B�b1�K�DV_�֋�Ч*��e%���7�7��(5gO� E�T�KP�~T�-,	��
����t�C��P6Z0K1n����F�]{j���d:�2@,��*�Z(T�>'?�Hײlϣd:�5���M5�h������Kae���U��}��o��Ǜ	���s�H��),�D�%9�磻��+��u��rԊ�lpk��� ��"�>�pG�VϬ۳�]|��k�hgN؇,�
�7}L�Tѷ\��'��F��[P}���y�M)��N�̙OёI󋥌J�maCS��g'd�	Vэ��mr�h0�&�����F\#��/yǦxf������R��8�v�.G�ye�;Nt�r��N��R)��gb�/��i��Gs�ȮSA�q^l���:���K��.�o�.ZX�c���2��OfpS�uY2J'&::}�,��
S�R�W����R�:!F�~�x-�����O&�P�ã�L�sA�lj{��(lL_��EV���ߊ���y#!K�o�bg��bZ"K3|_9`z�9����#k��R�u��b��	�����Y����s�+�����&�`��!���w�@TdR�����7�絍�Z�����S\^v��4>e�{;���kg��j��O��"L'v����Vfr�ڢ<����9��z0D�u�!���l�9_�J!:������f�{�7̛t��a�f��!D���'����ǁE1���/	*��2����c���OM|���g|����n�'�j��w�ͪJ���)�9A2�$q�kۈ�)y����]��3���k���V��C�\Ⱕ��XZ{rO�\��wЕ�o7|Z9�s�.L-��)����|q��
��Fa,tݑ�Dߌ}u�>�H�FW�4J,?�'�]��4���Ҩ�큦�=ֶ��!v�,�i��m{�d��$S#L솑�$���4�Aɶ�_|���mI\�'�@mѲ~<p8颿~R���?*8��ӹ/��W�HB�����2��(�T���M�!��H8w���6�g����8���a��;4>z��͚�%�st�o��-��@Q:�U�No/�Ȓ���j�"8T��!~����_3��_��d?`�K�ǃ@�t��T%J�vXp�k�I#ᵃ�������B�M��=�GT!����i��cd�����q�l�jA|h�*ȉY�?�{/Ș��i��H�'b�$K��a�ŷSv�3'O�]�B��E��On(lZ�Z�����.�)��ժ��U�,�U���rj:�*K
]0K�Q�-,>-Be=z�g>���^Q�J
�3�V�4�n�GB�����!�M������5��E�s�o�]`D�5[���Pe�*o���b���-/�Z�|�4�I���w܃���`[���sD%�� /�M���μ�z����4�NT�Tp>����ޙ�h��I+Te�ڜt�"^�E bd;�G���<��q"�k�U������?�Q�O��gƖ��I�"�<�߭��G:[���6�L��I�|&z}(B��_�nGR�R�Tǭ������o�B8��5X\��0��O���?Vt��f_�$1���=���*��F�=���^��{���a�����Z���&|���Q�&H	����Ӄ�g<�lϨ�{�b��C���x��!J��[�"�����p��dYܟ��B;?�4"�W�j����5�j�i�v㾅Ǜ6߫['�C��k)��s� �3=��D���F;�.p����d!���Ta5$ƣ�l4L>���똲��T���	7�G���Y[p�<Vl(���5N�Cs���zd��&C��Q�oe�tAx����D *�|�ɦ"���V�0T����Rb���=�0�>?:�hoɝ�z�G��
����Z�.ϝ�g_���(��j��O�ڶ��9�MdMqW	�g��uf�D����	��4�9Di�J n{kr^�1��4����k ��QQ��� 5�}��%f��������`x�o��`O��up����g�"@b���,��Lv'h'$��h�k�4_'?�I,~�T���� �̑3	��o�R`XER���2Q1
%��%�=���o�U+Gvߨ�F2Z��0��@�����	jh���A�Rl��o�_����Ѭ\%,��	5�%Op�!�^��^�Ug���L"(ߨ�:�T"��|r�p�Vq�֡�=:$�chq�B�k��M�����r��=������&=rG�q�	�hA���^�Ds�!��=2�]? �i���(5&�pz� ��"�b{Q�+]�¹�i���\5��9@곔iF�VO`R �P�Ԣ��&�������/�It�н�O��ݧ�b���G�n42����6��Ȭ�t�C�!)"�����@P��q��H�G�;�u�<�?�}:i1u��yg�EB���%�\ O��
��p���ʯ�<	���؀5�""O0��@G.v�]��,Wd�jT�;�B�����?���+�l�kA����Y��YN�zn��ՙR������ ��}g�y.=թ�WK�o��_��o��:eqb���yy%a��;�ây=61��W_W{+��g3N-�����jM�)�63��~a萟-�.�4EѱB^�_,:�F�Э5 hբ|d4�UW�6e��裧�	x�5�/�|g���q"; ���B�֑��ޢ�D�P��
������`�F������@�GH�.-�9B�w"�&1��X!�"M�=��=�Ml%��^Ίm> �`Wx����6�)H6zNO��Fh^�}5���q�'cr��'2��S�?�_ќ�NbZ�2���,�S�5b{}��!�a*��v�%-������(�
g5]�K�Ik��E�Zai�f�T�����	ҫ���?C�[�A����Ƿ���N�W�ؕh`�
R!����k)�
1d��Thp�*�,�:�ʔ!��Ė7����ɷ��:'����g��l��ZW="qU!+�1�c�jY��� �S
����⯃��=�Y%�%�H������ћ�ޭ6r/�A�(��Mf��ۺ�����K���e\�x���6mѹ���>�f8M����6����iͽ�x���\.��;�S���@3pq+���
{��oP?��˘�h㉖���j�(b3.��Y���\��4u��	Ek��n���g���b��n|?M+������a&�S�}F2��"P6{��|y��i�{ĞB�1�?���q �ĨW�|�~���Cgi�U��26���vgG�ɴV��R�O8'�o��^JF@��֩8_eC�V�ߓu�:��U�%U���!�34��EȦf��QG �9��N��Z7K{}ɜ�Vh���|-�ܟ�,K��;���*���7�oXn��b(�^9c;�HL�H�~K��P��K���P�i
c���_���<Z��Ez�9L�F&�5>��
�J�#�F�ޮL�L��A|K�����(F��k	��W	䇼��Oa PC&:Վ>��_�ԧ6v	n[r4^��o;Ai��tsp[�*���O��ᨯ3����s5T�CZ��)kO��q���k0��Q�j*�v��h���bo?
[���h����@��z�p�S^,ªϜԫ*����}��b��p������ ��?�'�K�4Z�ĕ"i�p)d�*^���G���>f<\ix�~C����7J@���>����/�[~;���-�1�V�,��0�~z�OD����%���{mE^v ����&UW���U�4�t���Y)���w S�+A�eƖJ��j`��s�s�-E��B�t3_��Im$�T�rG�=#����F3�>��~[�QE�4'�-
�;դ�e,rϔ��$T���ȯ��7�l�ѝ���2v�tQJ�C�E\2в�L��O;]�����J��I�n:�@��������3�����5h Y��Wp���}ټ����6�Vp9���;�Ol��k�\Yٚg�1���8�u����vu#ś�t�����IwO�Bt�h��JYe�}���2�g��]�܈*�R6R���B~aů��} ��P�̱
�u���b�{�3:M�����Wc�Z��w� �AG��#��4?q�l(ht.Q�!�_Y�x*��FpVZ�{`�5�/F@fM�It����g뗻ΤQ1G��$�G����?�D���_A{��_�sG�W=�TՄ���?^�ɔ3W�0����s�ym#����洷C�ɖ�	� g'��Lzz�.ˁ+~�&_T���~��F�{�c�*w��)Y!�?pX}<ӥ�Ǥu�{�BM,F�[�o!����>SіǢ8q����X�3(i�P{ޒ-�����U���:�+���Ӹ���Y����1���N����w5	ӽP|�b�!'���F��G.�cQU���u����鰊�*QL�_2��� p`+� �X`U���� �a�V���܋o���E�h��Zm<u��It�_��v۴��ψMDUS?�\R��1�����y8�Ӏ1O�[���F�H�C��Ѱ�@�������֓���:̀ ����Q?{��h�a����Āl��K#�i�o�l��^�ίj,�z<5���a�,�"@`3��b���6�N�I�q�G�����%�I�ھ���|��(�KB�i� �˴�ug���W�R��ّ@�S��'닼����"ʍ�0�A�=��9I�(���D�:�U�{�?�;��y�}�d�!��"Nb�i�(�iďC�N''� <6e�ݢ�#�yμ�S?ahBѓ�;	�K1`�c���h�f�h�Z�S�pg�� �дHt�k���s(�|�Ts��	��\S�$�Rz�K� d�w��i~:��A
��Ĵ���R�":�u\�Q����ݭ]#{fQ׆u:�T�h�c�I��3nE�œ�ޯr��S7��K�!X
 ��{�-Q&���:�����~&�������~������r��l �59i"�{���u�"y��`Ѩ�&���������"7Fh�p,�9�Gϴ��UG�{��1�xFB�GdL;[მ��S�ERXj͏�i�K�F���\����0�,�w.�Acj�=��`��s�e6�ت��%�2�m���U�}gm��KQ��/ϻs���@��MA
أWf��р��PjN��OY*F���n��1!KG��s�0�q�o�/����;nb��!�� ���U�7(��3aMѐ��m�7f�&�����~8=?l�����C�,�աGH��5��s�����Ijg۔*h���#��V��l��%�x%2�MIkN�� ѐp�ش/��V{(�fKOz��uX�*c��}�"�VK���G�x-��IQ���|��/dZ�>�h�̭
��49���E/�����š��X�bz�(��z�p�&-�Z,��]��[~��gf�4p-��i�4Jc=T�|���Nr�b�e�uTp��7/$��\�����a��Q|���)T�C(qp��VdMp��Jr�����^���;������[������Iք���+M
>�p&'����)�����p���K������(ozk�߲�����ճB+'3N�����Ҭ'�C�	ҵ�7뢝��?���Ļ����:�Ϊ�za�icǅ&3+=�f?�y&�V�Y^���#��s��g�K���w����S�]p�&�o��և�_(*wwN�/�F�F:XFXr�[$��o;9勾#�rLvy�C�i
e�>���Y��"U��U#���̾ױ��d��Μ��[���x+����@�@��� �������׍v;�Zu��&�����B�i��� �I���Ls��}YI��u�S��h�4�eхo�k�RX;�G�8�X�z746�H�{�F�X�&I���;�;�Z�� �G^P�r���է�飼��6*"�'�%X�fC\%��zh���q"�����m��,T�D����1\�	�{C��h�Ɛ�k�<��6m��ޝ�͌�	E�(SIs��Hs�����H9�Ѧ#�a�z�:�{�z��ƓJ�}k�I��=�rB�����)U��z<1 T�8�bH�׳�%��U��^옥̷��!�t54��� /�dB ��i(����3�E�ã����+�_����p2&�Vp����KV�3=+1v[t��5�ͻ�Znr}�� p% xObSt,v����p;�["��M7����<$���}���O���ʔ�4���/�2917ye[�P1�k^�>N��F�Q����T+��9��ߤ�H���Q�/�La?�UB�Nތ#�Lj��\ty���e�5W��i��P07j�D� )��e��F�7�����L\�ѽJ��r�je����VR*����{-c��6k-a	w�$7 9;.kT}% E"�4�y"�<7�0隴.���?b�5�9b�nS|D�Äӡ����x�������
J�At�C$����vc��-wGo��jn�_J�`Ud�p��3hP$�i.�A ��cg�%70J�vB=ٮY���?��u�����ߠ�ߏ��Y�R@�l"�|���q�׼v�`a�eH��|�n�Q}y��`�~�? ��,cC� ��5��1P]�R�Y��$K�b���.R��̇Te_c�=�(�v�%���N6���*���Tf�+홗�J~�HHtg7ϷN���@,HZ��n��<��H��Z�������v�������U[B�Cx�d��!K�����K��ݟK�dB�&s�zYC���>I����O���-�7"
7��k�0je=�G�%f�R��G�	'(��6ۉmٶՓ#b���l������aT��6���c���[�d�%GJ �j�<=:Ke$���5�-IDm���@l�����D���8ĳ-�Y�0>��gc� N�MS�=0��6������^�*X�</Ñ�xI��E\W��Jz=`��ls�����[�o5*�c[n WQ"k�G�$>�2�������z̟o������������`ݾk#B���3s�q.�Wh/��k�Io�\r����i�j����ښ�9�����(.g�Bdq���A@�BVL�FfW9�"�5�(�[��8�V���8�)_�����ۚl�
�!q�JF�Q�b2^�&� [�_��B�d����`ʛ�s�����"R��$��n��B�7��<:m��T>;�b#/�Mlq���s��?���d��o�Ѕi���C.����+5N��@'ёіz�i�sC���K���n�=�mo/ևW�H�L��)ud82U�4��K"ZE������zC�� q��:[��N���<m�Kq@�c�V�����dK-�N*C2֧&�^����g�Sq����0µ-=��kv>�S�`ρK��O0��W�Q�v����e�� ��Q��rR8Ț���zƅ,������o%���!��qI�ҌlPh�~����5���.�=��zS2��/��o��$�bL&����QZ�:�4��/i�S ���W�d�q�B��HN/��-Lv��ݤ�a��5Z��y�i���+xt���S��gW$&�@��zV�3���Ay�I�ص��;d��Y����a�:p�R|��~_�G�4�^�ڨ��5�4w	�Q����1zu<�Ν~V擩�x���?��+�sv���*�]���g���u�z�����C5:�(P�]�g�W>BP��%3�����LG.'oC؊L�d�<��-��t���@Z��x���f���/g��A���kY6``S�!�o���>�@�R(���Z���w��[ѥF�*X39�Hl<Emjt4܉�,i����A�S�n���3�h���ߖ��1��`(&��ȗQ�F�m��;�Ӡ��-Ϯ�:�/-��;^y�#�C�(_�U����G@`����@�h_�y�bC��v�ʈ���yX7�+_��Ľ�2#9k[9d�h�<x>;�M��:>���
B§�\�T\��:��T�����2�$�n��|�9��ϛ�K�B׸��e$�1K�'n�(7
��>E|�@��\��b��l�":V�^�rJ�_׹+�59�������ʉw�������Ԏ��+�*�sR�C~��{��^��A4���9��.]ѣ�D�)�⠬�fw�Ú��c�.�@�t:���'jZ3��j�Κ	�=�pYZ?k��e�Ѣ� &B�=�f���h�X��8Ȕ����좸|8�=j[��%O�G�o����^���<���!���+��ZԆ"2 �UwNˤї�e������(��y^����8��YƱMK��Ng#��m/[29��0^=�<���L�[Ë)��6�(%!��{�16�q�u8��j����.�djP�x&nD��5�2Pt8��K$B<����$�N_�r�X�����h��>M��) �㎀"����Pa|8^�L�)R62N��n�6��s)x��?�� ��>�G� _`]dG��;oPOF�Yı3�H?��TB�@�j�ġMj����E��*��� �Vs���|!gRR	1k%=���Z}�q���%�Z�\aQQ�t��U�:{UT?�'�O��T�PX�yz5��.9��2&�E�E������)��O�"���x{�߃��i_)<���Z�-����f�%e�R��G��
Rp���tC
_�?����;���[l3�wq���=|��j.�2~��4\˖�- oOz���{��}�����+3yN�Z��3K�!6͋����W�,Lj9\����pҶ��Wl��o;�O}-A�r�>ԩb�ԕ���}M���Ĥ�	��\'�@Ѥ��U��B����nZʭ�I���f�}�� �0��s�|���1%�:��\��䂭�|���Qv���� �ԃ�q�\M׌��Wc��Y�|�I��o��g�E���+�+OuI��Y.��1`�&��ݿb+[��\/���CI������}OK�/��+��*��3A�5`)A.���1��S'�!�E�E :�|�S��V��4�O"���(��ѳd
T��X��t���ze���-�F���6hc���i>tb�ҷ�*��n�˜�i�q�|w§?�������?���Ы�����U� �Zf��{��X��F:��ّ��P8D�QvL}��8�=�U���ڀ��_&�K��cDd(L܊]�Kz���MF4��ĵ��zT�ǘ�o�>"���]vC�lw� ��)~֡�a����OZb��eu�BW���'X�D���uO���r�1<^@��>g�ˢC����R����%��y���-��I�s�f�
���N�y	x�������p�1b�����!vW!��
���i�YEi���I�R1�����K\�rGi�yTIV�L�ik��dv_ѳVч���Dzt3k?����8�?Ιb�#o�x�W����c���>�[+w�_=�H��V"���"�Y$5��BB�IN1[`@�fU��3����uIL��8�tw��F(mQ�<n�c�6���Ɍ���$���)/��1�Т���""��pFi�����QB*/�ѐ#����CAd~�Mz��"�ǃ�	37sH��y�p���E�����t\�έ�¾�G!�;>D�C���0���O_��O�S�fQ�)|���GQA�a~��d�q0L�sp��ڮ�r'�O�:�"���"N��~ ���O��M��}�;�H>%���(xG��ȸ���Q�>����@�ů�K�G����vdڒs��ב%U�A�>�&�ɠ^͍:�����,;cgTK�	�l���յ�N䯀�/+vhS]�lx!����)�s���҉�R��p���N��$>xe��N5���Bm�Pa#�	���B���e̓s�����\�ls�NFQ��w|{N�!z)#�%r�#����̌�H��ɮ̍�լ�������b
��Y�n��������f����b�>���˶�-��d�����O��2��\ћ�V��g�+4	!(4�}Z�O?%����E�Cv�VIך�p'Η�JhLf~���9r�E��4'��pZk��'�N貟vb���W�*��>.���Q4n��h�M�ܝHQEcyvm�1�,%�&ț��	\ۿزtN<
��j��-��በp7{|v��"j
ʎ�)�W��/e*��Tr>g�:���|�� 3�4��A��P`�g���vG�Y��ז��FA�"K��H��8�t7d}5Y�B4�L��D��a91᝝S�dQ���[�V�z�{{1=]ŉ'��.�a$�����8w�dX������-�U�/c�w��c>�5Bە~%��'�z�Q`.��b,��F����F��1% b�4sI�=a
6�s���0�Lt���QGhv����6�܁��	v�p##^G����8&Vתи������[�)��h�/B�&��b}ΌD��mu�Um��A$��7:1�����U�a.�)��S ��ő�E���<�~m��Q�*զ��A���A49'�zK��T�|5q���M����;B+�o�͂�8+P�2p�9tcYg,��4ٜ��_���$%�ža�p����m0,��`pw��Q!(�AMH�O�k�e�fs�:��t�8I��8H��QB�DHpJ~q7����)V0]�yJ���L��?�+��z�����E��I �
V,��es�2a�@��&�}�8�|��x�;v-���Q	o_�֙��Sg�������l�vr���1V��n;�Bb����g8r�FHSڶ��2pxT�ogt�o� ʆ��ō*���ZG��}�b�޴�	�_�ްj�|"���T���X�#���O��Ԅ0�#ZU���!�w�{,K����x���i�i3&��cp��!��&� s��~����do�z�����3��1y�zʑn1g<�NG��w�}�OT8AQ��sB�4f�� �}�Vف�2��{<��*-i���7+�qǴѳC2�R���r��1t��m�[�=���nf)��_\_�t�����A;��9S�[[�"˒�t�<�OX�)��l���|/TA��f��mW���+Ƞ!�-B۸���-��^Eۏi�4	��>΄i�ݕ�r/l�� �o��K��. q,��b�
&�����,��q�on�:iv3��	HJ�fV���!QlV&F{�UU$��t��{p��k����� :/���y.�	k�Ok"�i9U����f��-��ƙ�l�Ľ\ԕ�i��/���@�� hE��qM�ަ9$ݨ�R��Q�q�	��.j�|#.%��c*�� '����p������1)��7Ɵ�D���1���e��(����s"�ƧF;F&'�&����F�����.� 7��X��K���g0�������Q"��q6|������K)�׬��y�@)�?����JpW��,�p[��/A�{	f�ͪ��
�f-%�1s���C+ׅ��?w���p=�&rFp����}.U��L�8��[���`�!"8��X�H�/].����P\�{~AvLx�/5�8�/s�j��0�g�:zl{���BoO�k�Y��DJ~C�4�'���WX}���Qh_��ߗe�M���J�H��~�W���	7[3IS�����_��Y����!�₭O����v#���Ԏ�5������L��I�#e,s��TǕ$��j+�WǎC�^�<Z/����} )I�)ԏ��
�2�g�Ԙ���9�߃>F�.X���Y��=V��K�C�:γ���F[1�����6�?E�O�W#�j�)�VK�����8��b��v��ś�_�f.��E'T�*���x
����d��빿�m3����|q
<�V;>�����P�2��S��>2�M�Q~:B[�t��"��!0��/�3� $��?�W�x����;�����f�K@p�t�@[�y���FE����Q���onͻ"d�,g/��S^ �R�;ۮ2r�Mѡ�������EN���B������(ǯ�i5�O��=�s�A�A�.,RO_&7�f�k)�9TDw�M��~�g|nhO�)8��M�w���#K�Q���3<���&X��e�G:��mH���M�H���7�h����:��i��x�V��ꡨ[�o�����G`ަZ+ i����UP[�[���B�tm���7H��v�m��ʐ�s�w�a��Ɠ�����m�5y� E�!N|�k�dO�{ƻӵ���~C"b!��A䍛���w�\��ۚc �6>�BF�%�My	R�S�*�בS��&q9;暳��u��sj+)p��"8�Hs����Խ���X�z>�Ck5(ae�2��E2&QQ?U��*�U�!:�6�Z�:!�� �kT2[8���Hd�}�y��>"2(ӡ2;�Ž�)�YĴ��\�/k���R�}@&��
���S�)T�OWQ|��s.+��x�V��4۸�u����E�����MI ����I�N���f;��ē��8Nj����,�	%9јe��t���0�K\��#�u��΍�(�8'�8��q�>�^p7���m�%� � ?2}l�tkV�s·���g����:�c���;���L�?��iE ^�'� '�mkھCF��rtZ����}�$��3�rmx)�|Om�ݠ�oym6İ�4��Ô� ���`��TaԆNd*h�,4��L�s9W�'���_�y��Z�bk�F�B|�GB��yi ��*r[�LQ�S��w��m����o5�;L'p絙>��L�,!�9U�#�Xk�%�
� |>ڟ@{�v�k�����xP{�!�%߱��\����g��GW���1���)�Z��d�5#F�c,x`B��qy?Y�oJ�A�WC#W�n�CĤfg��AB��(�3�%�{�}a��\�5�g+S�b���htx��ZB���8���R��T�cZ�0���a/G�>Kud�l=��uo�$k{���3.!�;�VR�1��(k��Yт���$�Ma�^�p�hm�҄�"�r)S�6� <�[�&w-,wn)\0����	��C�VP���be�C�$p�6wo"�7.4���������D�	�mع7V�7�8�	��eW����3�\�߮����dϹÁA�P$�F�6�H��T�U���a�΃}��
��Y]�C���~�E�8W������Ѕ5}`;a�D�g���z�'⻼�3��Kk���*� N��