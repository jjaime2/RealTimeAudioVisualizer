-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DVGZNcEX2PjGLwdENvF0pT6OyZfZ9Rzc5sqbFi6jfJwt7LvV6DIKMB1e1j1nyBupj3Eo0NGeBGi8
jjzag+7JgVdjkie7xE8hgGI1g4cDzwazvz06odoW5QupyQc/9I34p/pNYj+xPPg56ZWgXESxKJ71
7qqfMavn/LWAzbI8AJIclYL8IEUErreasGJmaJt5cdGTW8SRJmTqfAdy37+F5vtrb15n1eH7FWds
ANM/fombFW1Nvr/TCpEPZDv329Ip4i1MBC98h7ykUszMy7VYmFGbP7JL+gBGepFbLAuc7avpXxFb
p3R5zuwb9jHLIQZ/fYDdmOspjWLHw36b1xOu1w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20256)
`protect data_block
HEukTSJOEjeWGuGz4AJXAXiz0cs0vsZWI3CRBhe6eOKNkOEWZge1bDcjHcWoNoOuXt84IB2pOhMv
EAdM7ynmKELcMMVIW303xOu8LBxdrh9l636QiAyCxdS2Oo/1+HNnSQutpBp6g9xT4OmtJPNmvkTx
DCfFAEucI56u/hvOCDi7KLkXC/7smX+Fq0eMobPnfKmXfw56fWaquHCXvygtzp06eImQnzX65BCy
ub7Mef3UaIkk2LyryeVEhYyc7/5u6rkDcQeTE9FEqjJea7ogidepIDnDglA8pmSOlCvEOcbNECh7
TMkk6ZtZP/R5nZRIgLCs8jR5iC9tYCOo+qgOuVbpjOISlhiS9Vuq8gVtgcfV0rGYp4KJlovyNc+E
cDSjJRHgThb9hD1byu23QtnUsnNMZ/Pe2CZm1ZQst1LeBTSYp0gmdREj6Tdo+TXYEWBNZoCaYx9p
+zcNyBVcGdSUNtQzof8ll7lKkPp7XkUG3rFuxeQ4pnSJaYrs6LNSmmT78NHPUoSttKuReYYBDafu
ErP3EFWVTXzFsO6V2E+1isNxZ0S+6ke69k67xO90/xn4WWInK6xD9iyex2ulRjW9I9zWErymSP3n
lgO5+0f3jj38hl+5JPYmZLEaN1VUo+syQXhVu/NyAq4fMQ/h6dN8nClcxJpAfZxKFHI4RYOs2Hg7
gkK+WusrROt5xnpIdMC3njTFLqxcRS2wuCf3fu4QLT7DRt8f6zjfpRcxMuEyo/n0HdXAu80Ye+fL
B/ENt1oi/aritVMOWXy77WclC+vTINJ4xttt76Yam/kvJaV2G/X2shgzvjNfkhzFM9uk3C0IDTYZ
sHKzQ85zwqG0V6Di4xQQlNWmgJpdwv4+/izUiVnKkDKWLRvjPjnMmN2iMG3ro6vZEhW8rws4J68L
ax0R4e3epW3khCj1/JEapDLoq40o/bYHeCeZAX2Omo0DVQEIpFtEnCZTzbeTqZH928M6RZlWqqmG
SBa1eJfYynmFoK19nvHebFHNXpFsRESvmPF0bGlQ04NKfROwKvoDbZviTYHg1hHto4RLIZ/dxbEp
NHLVwBKoDTI/hEOH+1RaNY0rkVabkjqNz00WqviCM6ZNV46+3BFkGZDcu32eeS4RUei9k+P5MuEw
L26BPUvGo0tcgUNvMsXbt+c7JmV22F2XjWewDcMLIpQrrd8S9UlOBkiniOpLjFu/naNKiEw9PK4y
cvV1X4h5Z58lGh675dqoUzA6Ua9WfSQUaiGCbhVkrF+2HB+x4qpvSTEysc6vwLB12w9I2tT281B9
0vGZgTKipvy30zVIkph0eb5zRxO+x8AB6NEyZEk+2WO54HMmrVJmMgpqkWifHN1r430/LfXs5qQo
eB5e5JXmdRhiPT9+TG5if+/KxW5WGMW54uPd2RbJO7Z30gwhaOSJUxjjgVxSZQGr8NlkK6cGdTHC
uC1Ft7DhieEhqRpdYRIbEEOjWE/klHDzZhthjQMltm8s0+EGIACok5Mi7NuaMjo2UMyApnwpv8He
XuSoTcp7k3G23yK5kOPDqX2lcC1sx0uSZw3ASbGm5fEzI+GWHj3oPBQvqXp4XiODkxtPaGbmQDjM
+4hugpW4NbWOJBgaFcSBGHxUQUM8VA0OBNFNBhh4wxhtwCEld2sSUlacFBawBOFlLYa6l52JCBd7
PFBIAUwZO36fTwRpEpaptZrTOaVAvaCg9mRbDtB5Ni9LxrpxI6nk/8303z5CbgWLsQ7fV+E9yRzh
TWPexIGuiFUDiYqGmDKbvZbHyDsGrvyQZJNu25cvRHDXWyzXN3JZGgHhWNQliZlnYCVJmyaUOnaj
IvfidWqhqepLfwYvm3+KR8yyv8/0Llj1ThddUANTMHjY/sWFHTdJayU5N5kercUFQq4xxLJBInix
93kB3SlJbiQxBOGDK5WJCOuu69/q9E/pRGgqdBiu3eNgKDtpgm/SygSrz4kW+2eqg42w9q3s0qoA
02RimJR2qInF1ZQixO3pNjlzMnZ7+pcbweah5ofWKqMkxxldq68Ol5xHrz9RHvTTFYUnRTTBGc/p
y7IOUSVdaoODL91cK2ODkYqJSWAbDY9VL0WdKUa/hy/CW8rHQ6ec8LsMuOlYhJWO8qpsyUew2v2q
U7FQ92ktzXCJAHcDtdrdSc6PpuDxYUNca9n2xXLpDRT+IYHmNWaVsOEfNXMc2jtlsmntuypdnZng
xjXI6thJDs+R1zd9KKG8UJJ9WxMz0zCOqknRf9ZPSm7OmzZtQtRuS19H91wYmTYxZzild+2vqcsG
tCzKGNCselsTGUzkUz6S7DtUR572I/fF/rvmLEywxkE0FtwRw9UDsZskmFUDZqxoK3Kv24tS24XR
eeeZSkS34PP9R6KtqReq6lmyhX4W9mNtTsk8Vn9dX4LWxcgf4RXND9oe2oBa4rvhSUUO/edPkAXQ
Nb0JbtFVKKoqwHJIQY090uaJZoXyGkPRbAoN7dZZ9Fo7YOpoF92OOiMX9gKOIqCrxlFY7tscFdPV
r+lp5EtzDnM9PHyGoDzLq2fgKLM7drx2yZXx4kEpSrcfhecWY2ALf8loQZ3zXv5FwSiywFY0bWXF
oETNgW4vjZMpGmvd7QMsUJJD1F3W6FGFHTOHTNYjKXKkDtksv+uj7Kuz2NP6txZe54X7LA5A+ypF
2PBL0RQL4VX9fBIuXcTiDtTlTJmlwOGtB3FSxZBN9HXsw/a2JujP3R/r1MNfiKq71E/p12xA2WW3
cxK+63Nakdv6YHDmmUaTvwCdSohZUQPUcPZC4qTfLLaCLFrBMNNSlqwjQcqLCu1BCIxeq6wVqA4K
3PUvLvuIMEfa9cYUfOE7m7z4COU3MEShecUPqrp+7n0OOwmFjvL2h8dBxFfdrGeXBkZuzti627EO
SSVJorzUVtOeHDbxanFHTjlAwsQTFP5EUa/vHaCLssWNbY/xd9BgZv/ZiZEs7uJdFlCRogZEGgyO
mj15c63SCX1HWy4J1BOVNvGOKH3gqLeqD3JkAU/mnXy3NZkuzPmRLf7dsXTeca3eLiTje8lRtkGK
kQhHSSpWMdOlkxjGwZn+IWqm8R0jfNd3MgOuACM07roCjIGsjP/bk0wID0TEiE784MmbSm8D3EDy
9dS1JpqUbmbfbXeiee/YvuAU9luuOn5RBT3HPqaheRbXuCQAkJbTml/zQwZTiG81kJEhHQGAU25J
GrrVXIdRdkTFlgaYTXjjemTLpGIegKpCeoRWaPnqCNFoHv6hGmoiEfQ6yZlTQzvKFZFLxXygNWED
dlrwyukYzIQVVV1G5jMrSzye2+vdDFRwxCwsX2LymsLyYXMCGzHp4sfFDkJWn49GwevK1yIXTp+y
0rngNp+3N1FbJJwORJlix0ceO8ZBT/0FDQW60jKNiXDyLVWPGjEEIuMpTET9BjErJFbpCjdnK/WT
aMYhvXwyZdlcPdcuEJJHRhHDKoYOQJzznC71vz6WuFfoPuXzn4ko2tNV7xVztbVom4XTLRrNTGB2
boThywMs44+atU+BfYdxx/Bc7h9hrIDIDXaW6k1iMKJcr27MO6maNoLhegtzR9T3X0F7gmq8IV8C
7eeDWvKg78C4sm19aCs1x98y2jXBJSe0HiEtG4JOSt2paPCZaUrVb/XVY8/mzxEpCEdfozoV0dXz
c9ot44+V024SoYcaPPCUBSgbCcg5mCZEpR1bfXcYIRQXZcqIlHjJzwkgEnAxzCLfZKAtQUbJdaU1
2CKntuOmiv3/0K0YGVMH7ufI1LONpyTFhfmRs2AkU3AoL+imANx+9UE9VKcoywzKUFuAPqw52bLH
+2XUZjEO2ufmpugiT5pRjdbKb7FvNNU8lHL7LhvkX+MdQIH0G+MtlybXSB2MFNdo1mVp7FWqEmEC
S9srosoT79jJqCDisBXuJXvipH555XSJ/7EVZ70ATIficHzRMLlg1W8+SulwAIZMsPFoJordLxJD
Ts0G1V/OE2BRQyB9odmKm9jI2jAj2i9iKc9CXzxA3BoX/WzSKKtJ4lqyIaFBECi6zZD4heZ6lPG7
D45Ea4qCrBLpTfudGWqflOh/YAAWacwCU/vKoZMVZOg7cny+0LGPtcTeitMuwA8DiyXoZ7TX8VCT
t/hd+8qqQPAcHMY893B8AJll6mMbXIRihKfMeIufLf3OmCmLmBmPM7h+Bd3zhrwr/TB/dsYwCQFK
TJNLL2ky7Y9Q92Tx8ZfWXRPI8jceGtgxCQNkf/LGim3naYftHMlnvD7czlw2ZJRWhUDb41RT9/OI
FLpr5V0jhUngEk2PRvQW1QlpZqgxxt2jz2JP8nOz1/VY4d9NPI1qKti36atwP6lbMcRFR3R5rABR
9lEHvtLqK0rahiWEKHw3XAQVM0jkML81L6OLQ1KjExkpaiUAtJo8XwiNyE6GGEEl5r0STBlWVGwJ
vJc77s6Ay9zsZ/KPV+GvjyGLQcwRQvaxoOo3ry2tcdFEeNiYvmbOrJ3aLs8tmnId2j73Wo2xU89G
fCB34VbzOMHpdClPYxsCLTN/AWBLVp7967GL+4k4k8BK27fCfAdTqEzSACc3Ftb90PfF0r7C2ZEj
0z7QP87XFkn8ZoCoCieqESh6tXdfEGbVMOsetIOr5tSuDkGOl5rVNnYYk/SusMokD/D/uQ/MJxCt
k5UyD+SJiBkBuc9MOlsG9pRByikds7icJPYcD/sx1xb/QhDxegdR+02mRRHBXjKHnDBsd/BsqSEd
AanUlZqAdiJK+Iy04hE0omy6FdrNI1BYxc1SHv2+yc9x65PzquqwRhutyBD/gi7GPrmPt8bskz5t
CQn8d4mbMsxYX6ouCk9mZp4/5Fu/1fpjZnnwT5m3W7WQevaq4l6d6jBc8f4VQ/vB5wxxX/Zt5T+1
EaJYCgkTGOWHpxZDruUHRDNHj1zuaQFKbpOTeoHldeLw5rMaEZwfAy/8hmwup6Je2OtHXI1rTw/Y
8zE7h1yrpoyyo7T6C9PHq8s7Uugpmv8d9YyEllazVwdj80oNyKzs3955B+BmCncqs/DD6ZrsGtiJ
Keow9xAcJUhSLZeNlbTSTXGEugdj3IpgfZcayxH0ogyi+d77Qfu7ifHrObACmSa0URzg6WVqKeSq
NBOMAj1Fd7mKzzIl9R3cICEEMVAdPsRzNZBc7GDwimdMKVmbqfU7h9vr3mIai01+AP8k05jkaGO6
oiruk6kYWHaxtUqJGo/bEG6aRakX/NmrRY/VURPwRRhgeJgrKbDLFk7jiQAObG5lMD/GuqiNmE0b
uCBX8gT1tKNX/tL4h4UfQM2enE+83YRcR3bGg1OP0hQXPuiGMK/JNjy2qbxVy+nvreWqyTbJTo4Z
LMCL+Z6EOnXmFOPE3CTtrLn/lJIO2Q0aYLMgN35Wu3iMeehI4+UeiIam2S21Gg1yGqjoieMLhgpJ
FrHnl52D3vjFif7EZs8h7Vgo99pm2cZ90aQK5u4rH6//zvx9ybTz6TTTfM79jRGWqrA8vz6XNrcS
DJvfl3v/eT0qzev88T6353s/Ic5ejq0VgLetASISNJdxiuKmaE3x8jDOOM/6PTlL7/xpWVBDUJe5
GiXzEvd9CnPFGbUbIy9vos4MXsF8QWwsNGgffp2gI6uwCFgN5NRAG05aPa647xPrppIHp/BnB/J5
2jBrTLe0gIjKVjKZbnqpPQJoRrDdzlnKlVgYB3mKgb4zQVEvm08NN/M9uosxY7lfhDB3Wx3QeXHM
LhZYDnNNWJq8Zsk7VIks9aTg09VVXaQZp4GB9MbbAR3tUKQKypwMjN+5h7//AoTVbBFJJ1+2ZUa/
PHK/EYMpCzQZ6zue9f5Oju8E2agszlpncDnLUPH83j3TaSOwgKOZfq7+8pTg56pRv8YTf885KWr4
uGn5tTGl1//8y+sn3s2ks2hU16Ch0lNmENWVqzU6ZklB3TVcTRqCHAeFVru98Viedjiri0Z85xCj
A++ZOCi3q3JBcBEg2xtavul99+nuDuEGsCsq7GOqjGcCpFvVDpJn06l8DkeVxJG7jvGrmCndALuy
a3mvbatSrQq63AswoO0coKP/yzSQJL3l7Fol+nATv50hOC1Sr5pySB23QkEmlLBmx1gnWfUQ+9nB
N1mbI/bMoYbSNx7gdCG6Dhz1Bket38sKqrbNBBvQbgpNmvdUoV02x5gEUHvoJWaGwXWjj8ZPR6ng
mXd2KsjGt+RZDn7uhS6uAcAFkZORlIcmGZCXiMZXoEP0zAxKMT8jHMmpNgVAx3cFRGkuW7Pkm+yE
XWdR4hvszLatG7kfmhXto8VrquP7R1dIqChWOw9wJqa/3kQvL3RCo1FpoaHGXaoMPI+G8TV9i/fo
d1DtatH9nGSnops6Xrl62pN0+pwSWUb7VAaY4kLpjdVDhiTWy0io3B4QdJjAmlzwvTVCkr8L61va
Lhl0DUTLzm4goxMEgAw6+98fY63Q4gVcovpEfx6rTiOJjEdqlpVeHPa0jQWChNViz/pE7ca00sG4
2o0cTywqi1T+3ClAC951pFG1nOntN1DRKn7VMvwaR6GVnl/2XP5PFaMCJSaqQ9Kt+qZ8OYISgL4m
L/J/87K2sjdpHWHEuimylyr7+S38joWcjjL9pVswoqRADJ6THpkjRlHC++9plucDYqCs3BfWv0as
8J8pGkzq4jxJw1d1PxAnb9m9f69v79rziL+SMgCDJ53D8/HnUc963w23hMCXZRImgQfr4O33oUcG
lsTyYBwjg4Ciei4n2fqpa18yBnUb2uKa1AiFRf8af4Ix8UTK9hzEEAZAOWOAKXxyTwDIwA5PY+D7
0zZm0of0NT2ZgwScts5x+mFuDY2tAYvpmdLiNudMnv81EOBTjBZGy6FJM4Bd+xM4XdphGppmmFkK
VHKluOLVNnHGFtbEeiJY2fiH26riW1WGeYM4lmZPNQ8ZCdB/P9WfbafU1DOQVz42QaeDJY8cEgsW
ppW3wlP4shdJi2b6spbTQO3F/6wkMF1XFSc9b2RCu9fwnGo8UeoYZ7huJ8OLppXS6p9M440kB54R
nvwGjoHoasIiMzyP0wwZw2gCAT54qks/n3QDavLK2K0jvHWauOyFgdBopYydNU/pVSkbkzGmaaaM
bGGT8ldch4S4T1HLdImeWcaxluKx7SWfa4vNQ6uMypuP5OuZI2jkNxPx4Ux0LuQOYEqGTYTFyeCW
fSAkZRJhjE/BNxBnSoN318/sdMOl9HElWqCs1aCmbfPVP2p/hYWFTXOKEFeHgoOwV1n3Fn++C6fV
a+gDQz9wdbTcwL6fqHc+HavsPRmh8PDCnSJCxbn86nKASLfRyRhsl/C0iWTv4Ia7JxG3U7PIZk5D
aJZa1f4y4xkA2ZcXnjHLc0fs7xZzbPiGn73f/NEakeBm+QbQCJGNz9GPB5KDLRguTsVrxGCGr46a
pCzKMUGEALAJ7BzmZBhQE3vdn20aAIred7LPIfJE8KupSbuDxctHqursefxVW9n08APXnb6owfLN
S7NKDEpByzfcTyuSrjaAazcJeyBbiGoCkEOct3FlJPArvA29B67GnoaJdLPJUAgoUflQb8hpi0xq
W8Rf4JLPvWbq1lgfB0/eKFGnpRksC/6yCtEOM6oHje3yHUjLY9O6BfU9HKZObp65Tqct8fz5AYD3
vAhHC8Eb5lOjUFMa74YnC70e7aWzFetArtSgumWmhbj70UPYmGmO+8dYPAarIcDbkiMMVskEpLXO
zL1TZuBDXa97IT3BnLzewwWEJJX4EKRuYKDVx3Otog2okboXHWtQhVDZXqRAvEQxP6SgumrtCE02
Ff0qU/tHzomdK1ehpvJC/mTM6iz20uS9FX36cFzC0zIRHG+/sRUm3BdNBgh5gCQPQK8/eJx2l1yy
khR11DumBj92CfnKz0+QzK5+zOgVnAODjFvgcVXaJxMqzGe+fP/C4V8/iTh7QVq4y44bwJn7lfE/
nYICU4AtEEx2vDFl1AqC9oPixJJRnBMdzuJQZbt0vMt6eaEGNKOcL7HVdtsWIQVZxQPYlOSy8DfD
CiNRnbeuyRkD6HGzyYrDSGuvFVjkWOdTLeU8lpVX5qGefCtG/lXnma72W67eKn8oeFxryVAsV5sw
VmZ6w/q0qgf0uddrAEzcj1kpqTjKtoNi/eSL12Pwwff44fprIbN7VeTwNJOibI7jn/CAk3nKUWyl
l0xEmsN3Qx8SyIyTIWnPwq3AGUefZQ+WtBED6Ga8/RXJi8vyETtO8QB8EBJDwU30/1pSSdqwVJ2v
ikPCgm0fT1cRio3E1F3zaVZKpPP/rZ/a9cCUqNtSYMwkEOSV5UheA5jr4bbYPxCRXa9JF0m3ZlFB
mHXRvbrA63AfWsgQXO9APggYwniDqvh6+eEInkV5sie2SG54dNuSOzD2n1QKjfyRusB3adO/C9a5
y2ysDhem0uW6uKZVuLGFvfspygTy/pTNDfm/+OAdd13ddeNJo56xEdebRj7ZMkDD1C1C3aO8gMQ/
Nbp+EtI/gEOi8hAC7iPkhyXjmYoNlhmIVA1JiJRuAA0SQI+PMq8jHw3PmwHAS2zqc96o4UpjvvXw
18/bCH7CKhjL+kQ3S6xXzJG4U4BuDlmozoLWClyrVA/HqnFN5K+7x1BhsQUruXCTOyhqeUDlZBYA
jccVWY4pygwfqM9nz9z12aGQMslObHN+mhwf/3L+33t1/iJbnEQxjvCHfJ1l62QnSvY+L55WJ3hy
4sBxszl4pEyTn0ZMQZ+3SspohNb5oXgjEj+7JNtORaZip3Z7lIcige4XlPBv2WmwxB7khOuJRhpE
ldZM5Lz1BhRzRhoLQIXQi3ZT9XKnbZP04cG0Lfw7dtdnWbJ3AhmSWuOst0qmzV3k7qNrvX5SA2gn
VYPybuPDGr4oZVBcS8MxFh9UIaQqPMZI3c0M9uoTNTLwXbat1j2Y6SPgbxHoQFWUSMfyp38KAHdQ
TM39cgGgvKLR4vlyH9NFcX+pSOf0X7j8p8RscJ5huoatZ6ehvaKc0ZZgbgxqMruAkWtZ3RKYt775
HJW1dgLBlRHLFVFsisBMGzPDitHgCS6o8lmwGgGhKr0j/xrxk05LRIMTJegxFvJ0p47tRb6bHpXt
BZRWO5sG56EBlbKFl+WiPhl7boO5Fixt6Ln58iwIDffZsdZmOoAX4KS/2H96rcJ8IdM5kpffQiJP
/X9ZMVIbghWgGfyuAbf2F8cLFkHk5uJlLw9ABdTPLlO6s03E23MA9VKnL5rWwhKhFSqzRfugstxh
sJz+2rXmeAWdWJS6D/mi3mYjsm0nfQSptEYSN2FMOsF5gF3xmIiUz/u/IhIlt6iXMIq1N6aQ05yV
4pCZyWPv53L5ce7k2nFS9z8ywn7vI6PtowyX9xhwKabWsEfhvgpH7rTCnVPzBiNRZKfoLkTHEeaR
V67mPimWL3iww7uioI857LuBWrf/+Jdsrgx08mzjc20Mqw/EO6wb8SDI6zWqjJnLMH73WjowZJdL
Nd8DwWoogpeVWZdUqz2fj8+YZOjd6Z1V9lMTOr+t8V065nF6jFqbjT4O8mBLh2ToCtqe3qSbsXun
w1p6kzldaZiDjSJgP63/T/tUt10hzp0wxVjw/NMaE9i5+Y81bchVXtEKM7bHGHzBmRZALVBRN+kK
T2gmBinDLwczncBIxV36J0vWMQ/J2f3IV5Lassk/QlASyqvNb+k3w2W7yXV/j/WMmDq40kMyru6b
FfCNcczhmRGDFSm0PlIx1an7bFtEXRCYoEvgkt4jOzpzkQTsCPJM3fJ60xcTbMx5V9Ynq1DC4vsK
DW38EmW6IFAB2JP5LR8Dt77tfMEQtha7/d7TBN+FlAmJKKd45uJGakemqusBYlS2rS+O8q/TDFGx
gp8xYkMPLn5ebDyj+I4EBQEGEX7f/n3l9fIhg9e9YseHabGp7yvhD945iZGdY86GS8e9MJJGb2a5
vXk7W90zVkoANHQK2x16U+GgixH7ACTjffXiGW32X5YS+f9zJLYVLBGFdgr/69LR7D6ddqo7KoPb
DU5xIRRBzlEYnCQrC6XUAH07paCGNlpJBBBm82VecxhEZYrNKp5ersyddM0TUUzQ2F67a8v1jyhn
++OH9RCnOPjLhEyTm8hziMvvHuOZOmQsz1+zieDTrXMNDCPyDwmowOeZQ71m7OADI1oVH3UZKT5G
O+nB2L5IQw1tUNItiZaXw82TY9KMWm9oXume81GldtpAovzZfzkWyzMlJbcC6HOchV949UwD1hyy
V63lrwvSqrm3OLpylU4QhyiX8ugSwjnw4RMxBhnK764/2rt1fcCdHlbBW9cvqvDasV5xYzhH1vks
BLz6LsTkrtNqvUKYV4Z0B92azce2sd9bjb0Y11P6/nRvc8unfuymrzHWwpe6fXoga3s7TUz7zLvT
9X5GNl3eKlNL0LkGGIrAFXIdRBKyItbCsp9z9/I/y7yVRc8sFddTriCAQAcVoICcU7TUFg5Kxt+D
XR2Byuo/Z0jtSr+U5DbXnAiGQ3ZYIpgkXtqkhoKpI4ilMkJFXSEFbib7Yy9JGE37S7jghY5JNHp0
n0DlYLm8CXp/UC57ZTjdifNeTouNbrznWAE9yaNAJACogGneKPgQ3wr2amC5tJJorh2mcE6CyrbD
lPCUZNSImyJm6mr8HmRgceRamGMXTHVcyx0n3JSOrQ/7TNYO2ce07ccFsqieaf6LfI+JRgq1etRU
+fikuZupXSDuMmD5cFTrb5Us4dkJOzJCcmQLNoxaXXn2Nrmrammydg23/9x7Uemliu2sUUpJ56c5
4IhHI78JxXs7cPdZ4Q8eLyKy0w+kpST1l3Cz91qo/a0OrUQCxKwFOPrus8GeRU47ggCOGYSWGS2Z
BMfw8vAQ/KJhlKLKUqWBEE8zbKueYEML3RVnASu/rCsKOj4FHpVLJVQ1Z7krMTSguME1EgVGzuAt
55nESd2r/xKf5TvLS2l0HkbBKWGhb5ie6JCg0LmilnH5BOv0yeTQ8iS8tc/odg9IKoyM0NS4hCCk
3wMLbdlkbIS5goy1zHmOC7LChnHPrFFW+lnB4Pw6F1QandhFKmt6C+96WwM7EJEzc6cG0++aGk+v
8zTCJB7nIXexEH0w3Yuyij6cLa01bc4MbtiRFggJzURp3QKHp39o3FkToAQbmNXj56kdThzjLRwk
+ZJYEXEDgUB4d67CetZYBY8CKewzBp9k6IXaJiSTxHI2FFAIORIvEmJ6tUgH9+/Go2ief3rXD/pA
ky6QSb8aY6y/twS+hR8ggtTGhXd+uI6CX07VBT1W5Rcy0tK/Hq6wc3KoxoJHlFMqrE5ZvlyXzHkH
2TfkFn6zUBTOIGCgPeSIq6n5QCeWG2Opd9cLFkO4rphKL08JqSeUvI03+DsmpShGEQqOxQ/R8zF6
cJkw9wmvFUCch5PtjtSpBSYj4oRsPxytQQjJWRTvhk2EDLHn3cUjfZnDqAeOzBi4HoqX+tQR2Svr
oQYDkdKAWYP1dDZwzxgVZpJjgcwoWzg2QkSKy4CvgJUCfsAZRZlLvzNDXY+qnd+AHDBojENmVSIz
zipSiT/eeMPpXi1RLw+Sq6/HImLpIAZhOx1jouVkeAFg8ju4xQtoEt0aASNi4VDj21nu+hqwT7lZ
ZKK7R2HKOZ93Hdo332ZmmK7sfLne1vyT05A7+F+I1gvZVZAVsUZy2sKee9jqLYQoeRwE/5iiMvIh
7offG8wsnorpk2gIfeQKJ0bN75Vk/dMIsuc9ovvPNDPvKOC2HRrDFrfsjwHYcSapPecqJ2hAanr5
nYMhqkuyUST218If0IYaLb5Vg6Zo1MNpr/l8zXrgsI4T+hjS+Q2ugm+nXKB/lEDSBE/FgvCtVEYt
yicXfkE7COfzFw2aw+6Vgxo9Mo0sWoV1HgU3mWE88TMzmIvIFZFvKMrnnpnqkueeSyjx/dnsilSg
CRcCIIwk/ntK7zHrl1QLFiS9meB90hT8+2XyDays4XZWZfoz4DnTxSwPo5Qkg+tJhELHAJQzFM+H
TogsuoMB5kMzbfziEdBW8LOUtSgH0MRus9BiFlOKjaFVb7a4Z2vAXmEtPd3ftbQDVsT7tvk9Swq0
pmSHB+o+mGhV8u8JlRtf8DmJuLvcgoKybSKXeeVZ+ZVoHa9aWt5UUJlsiC04idfV0jNi+ii+hIqf
/SCdsn0NB7FZnJA3oyR+rNXIF8iO1JDokHT6xn9zWqnk0xn3qiqt8vMDqBAtYIATaK/OwJzknOD2
P1gEtcU1s6OuHS5EmVZNyh+x+JjO+r5et6YhlgSqeJub1buFL2H8HdauNakgoXmcFfTtQenBeKUu
LqZmkOQhNNZzRGwNlSUVXgLBCNyQWDC06Y/o18v+2l5klkA59E2ANID2vniB3sdMSaUSWZEtxdfz
gi+NJxCOGVD7n0G4xGM+8nisJrc+sKbMjDHvSoLYJ6i9JIEV8RSsV9GXL+Z2NF6Y3OydecIk7wJS
xIc/hM4Nt7vyYWu2DwBW9xmBkqSGQBf8wD39dcrSVLUhOGSzg7lI9B0xNhtVjyZdKVdYFAnOmFC4
pxJltY7TH0LkK8k7aqSsGO8rt6cfBoWdzg1Kv3b7TsKH1Q1J9upqHCJOs/yvNlJsLBgXTmT0QSvb
fFy8E1ckCC7kXINjzgvsgeQVUILyZ1bHsCA6CcENTJFTyH3Bv2SskPzz18B8kKt08k92zRpLtLRM
trwQf/2GUqfStmehgOtidZlCaduAZR0YCl3awuNH6zlrVHv7xaGMG/p0KheO2SBQb4CTJURA6hG6
4jap1PO87iMs644Xy/JxJg4/8yv6nf28Iwmiy2HMfqHnPCw8HtpvYLctLQ4lTkLgZ7lja/PkQjjf
SsHMMytCLYTIiqUdw5gWJkM8tKBInPyYSxdG+MpInj1wQRsgISI2Swe14zREWcaCONZXAzO5RxnL
doyk1GMn8gyxIGOHSsZ1daG+Eb2cV91+yY606n89Jwk+tygb6cCfkElx0+krTwm2DQb3DVAsCTHd
ylSeGkZ7ZichJmdOqz2s9eSJJYyXZHPWo3xnKphyGC9QlSlHYs9fLk9i+XQmsegd/09pH6Idb1LQ
frkVPAJa+hT31fT3qWUQB5S/q/yZuyaU1dD0VzRAFOB7p+1Y1maV89KSosAMgHLbq3XXsDC/rFi+
499ksKVOEVUCuGA0VZp6+zOKfx7rLEsUh9Fy1YbdtTjxjj4L4ihh+O9jh1fLan7s+LywjD+yZER5
WM3dNXX6cz0COq1J5uV862myZwiA1DaCggRg0MybRKsXhPD/mi/kThLRtYB1WTAAGjLRcu+szXco
TgcaTmhAq0CGRekKc45hs4utd/mEGSdloJnk2OPHint7sB7TzYw8KyUk70W4xyE785W8sQ9PfcGV
8tC9Ackroko64a8Pye0HNPB2Zr+zg3HBLI1dtMP5JQM3RHXRhS59hTm8FwMP1HS8VThlhbBDa/Hq
2aXM7mOz4wjCPBBct2d8kqLxEGUym2QDvnJNTVJeEUkjlk+bDJA1A68CgK16RbFR2BBcmgl/tsqB
eP4xK4HLneAV6Kyi+s1g4bpuusZFZJ+TU61qu2OQM9p7dGoFsUaaug3IUTiv1t/+NgQBpinR5Yc1
WX3OlBASkg+vxwlljlnZIiYQqT9qNkXdx3JEOyk1CwGISM0321wvO2fv2RHUbq610VupvIl1uXWt
eO4bV2/7PAJO+ux+S/YKpICxiAYGWlIsQRgH0bn0NiOjt5vGf1qtVDi0nSwVChubID5kbK0qgmXI
VyUfWU6u1jwFofBE5hd4RB+tb+9ceVdE4EmM7mQemtL1+5GE9Q/thHC246JplyVjaE2Xl2Egz4Zk
pGzQovApwnvDIVA4CZlD7kZbd/92kEVKdd1styKWNlKDd1MystQHvDd+8RAWog66z0hhX3flytNy
sCRc7DyQNloQn/Ju8X+SxPWGYv4XJBY1SKD9nH6i/kKR0wje2eEsl4OgPsMC6efeDpHTGqf6L0Ob
Z9AeFU19dnaIMnZ4quAySLD+aYEsav2kW7Ji2aSjgPjNuSe+nfrv0cOTWPa5SQmCilGkjwGf6zT5
sXcoe4a6tk1NIWmce3BxxUEonZpiUuGkR0X4ypAdcbeKfxe8ZbTCbwdyVnBQDj9pnZHKKvFr4Hji
hnh2wCryf4p28to+xgCbj8ehA1g5KNG5JW5Rj711ik6nD9lLQaFC2d6/5LkZMVxOl0iFtscMz/Cx
ZX/grf6pWFC9K0yOOUTcEoLzzT1JlsZwJazTVPa7sQ+MOe/GxGqQFVl9/bxJnWNxdv8fGl1i5lJA
+kkrkzJ812mUGP6zToMHjcoJFd0Bo2RFrNcyrHK+xpRSzHNOBsqfkQ8sJJ/q9LxCsXPVKvX1GxQb
15aXQ4mHVLomxFrTkJfpXH2JbOxLBfgpdD/KV0jYTIKx68ZfmxFAzgut8mi66VE2Axoto2O0C5l3
fD7Lf41OOi1tfZZ+epWdwmMd3MI3GKCDqinH81lAI/M5IA/h6YH2TFgVV6cA6Z8p/me5aXAo+C1c
Ca+Nl0AIXnrU7o9c24gRhFLKJ+tkHmDngyuP2Z+JOTXkxKY57mZjOw4AZjn9+ik+TEnWRz69Ak/M
tXt4WWV1sV5nXrRig6uW/gTXBVliXAVCYqiKYgTLK5dUgO4OT2bDRhVZeZR1J4z1S/OloBTkHZpX
Z1lqgQSFc1pbR0MH7+KWV10ufNr7+WM288zYOmRA9Ft/++6bYg04Z4j15XqE1GeYuETfrcPlxhE2
NpwALfL1qe1+5JxxEC5Fn4bknvY8uIs0Da4HqxK9m2Lm5+n5FmIanC/7Cq1PfuBNk2NwMyUROJxi
uUdi16M2pPO8AwOyN4aFTcP3aVRE/KqUfhG16RgVxc0mVNS8yIhtCK0sVzySx2FpEtbUWR9ziy/N
clroVhg4uuS5lxArCQemViXSVY7g8LrnQrEzTrk2H78nNoFydrattImqDAyhQzi5zxx6ik+e71q8
2J9u8YfV2QljxRCcRJB0oBOXMfSF7Tc7dSWtIGpr1iYh3JOyOcdhQ/2bOJiJedTGCpp8andkXw9t
s25z987dT0dLsmac0XRO4VSd/K6rk1VDx5mlSI8t4D14wzGVmP/+d/URrO3F+LFAl5IgFtDQtIHs
IMklgQAUk2vyhC7vRN0ri/KQf/54pW+ik/0hu1j1X25DfCxHcwoMU035jTAvB0ml8KNSkxWlC6VU
ApR28rcndjZCNZxPLGnqSrcCwzNeuQP6F+LltJX8LfAahHRIyHGlW8M6W3pGf8OSb4bM8pc9WLsQ
1TyvJ/B1Tb7dyfJbxORFGKZjZPXf/jIL+Az8C72PXBnoaKGUD3E9k/8xbQHt26ngKAnYB5HCkM0s
yEiO8uE9co2WXK+NskyYkfKzPzK2XZJ3n6RjPYaP9ntk+Bq+IIavnhvtL7TzAZw/7U67G6R4YapL
RxFY6dkKXTiZdzQx5tHsfywSmSkiKLyuh2oRdd9hqINg7AIe24HLssLlFIUW3rmkr4Rt4GXRHBX4
xLLd+PeeO6by6N1M6iuvFY07EhUjlfQGQQlZRz29+kSqaIBYRLdyTgnQhJk14xe4Ji1Zk2M+raw2
/VbtY00COX3VxtgYvg61VplaNFCFmleflbSWReYDcPgFnjqFKsCcIhWHwEZn7s2HmqtxcGHwtAOu
ISPBiDnPwxMpihfIZZIUbpp3ECtQcap1ZXlxYbwWK/KtKh9EUSa8HooNa921KlsQSLbZKxBA7Vfu
4zszM8JgRB6sOLhb69+1Wf3Xu0riOKUrJ0scbZmHJS4LCTF1eNWlh2Cfs7N6mDR+091PXMi+jNJ5
mveHUakig67UI5F1G4FeMhSomMhD8/UxIzBQHaJ20HFsNaYf4MuyVweDTTSbyfL+pensdWvpRUJg
WSjRl4i70Pnhk9hVjUFAIEkH7dC4B25l/emD33yG7CxtrN3GWzybvFNypbXKIR8ETK3X07g2asq8
5aC8NxXInv6nrzDqXAgo7TwA7OwVpOQNbXZru1MGDOFVXDWcFg4lKEOkT14SZPfwiIeIp09TRt3b
TOZjqmRRGMP9VKlrpOsjHxvgaEQmR5zdRhV1YPFAEPIShlyQCDgX8350lDarvk/meHhVdwmAXJF7
YsHQrPvOI2l0jypwpvqGc5XEQmXkD7LO19UnKThgk4zO34aPU6zovuuIcPnR+smCLtjkCJMCLqrj
QkpnAUaPqyFBntNz1XHDP+XNk8pgtDT0SEI+IEGs06o4YK982SMiWZ+upGv6H5Ss4zHzgJEak7sd
0d6vlb9ZlGH+rDMC3oEKelM7aaw4ckMpyV5WGoVoSeelmrRf54xOyZH4UKF5M6oC7PJnAYM4xtL4
E0Mba0pM2fj90msirlspcC2Hbpb0abdZCpf6pFyPZyKjOOFpNkqWUwdjH7wn0NhR+moh+0AKfoI6
sHDEi4kKU+e6eMN5iX7wrPkqz6Xp+aCYdSSkZhDEEIbTy93ATn2RFg/nKea3wliAZ3hlkryEG3yF
tAMZ8dyoW8lWjhf7B+zxtfyvVwgdkjUwWybw27NtjbdS7O//EYBJzK2swoeQs8Aa0zeAeJDRa1M9
KtuL88Vj2yHGcAJI3vfCUPwIGGsdDJMYqp7/OOyN29F6rqyTK26tmBiqK+DHNZZNr4cokaH7TNhP
cvXNsrQW7NmoVHjYConf89ixBwMUKG4lab5l7LKk87t2pVje694Q8DF6dbLLT6wZD9qSPXCKbW5Z
VhgX9YXh1aoIjPyUfckScbDZHsVP9i2x/GfUcAyyZuygSAUXP2L+28g/pZK8lEPDzB/LJFWiQXqG
3Rbiaa4/dzQoBS+valFWICL8KLJ8pnYHKZ6+vKCGwioX3rkdvfzxAQNPOmQChUh1ZR/1AWJfayTO
dW2S4GiEuHqGIDZTBWbPH1pDP8+zwhIplXOiJG1qSzXkM6KY7RIZeGzt+58EvxUnzQD0P5dnPBzg
4hAQOHyQYxh0s8HSACHKpmouzn7ox6pqor+tymF4YjFSuCE7ns9AN5uYcOY0tpt3cKpJ/kqUf4tk
WdW1BQu1FIiZIbiix4utS0KzVDcrJvOKAMA4q1euFmqQ3ldU8dDWUg900EnofHGmnby9KTWHlyty
U0PQ9qeIoA+g504ps08ZaHyDp8mbOvoSRwBI/kBInN7IUaZVLCELmbsLiLVgpZfVrLe3dodnxQSq
ccP6PH1kjdxy+zOk0kUH92B6LMznyS8RHfFb1+w0dx1rPT/UKvvjpODmPsFyiX0Ayg3jIBKmVGVs
x6icQGwrr9DZpDaRJi+8tU75kF21jwqRJNVDgLg4NVaC6NthyFwSgaXwbmZZs/20vFg17vSxYStB
nXCOwZ2dkT9VXn1227ulU8mH4XtJb1+7hDZLC207t1OPJq7qJfMfaYtUYsRt3It8bhggenbervHl
wQq9/IRuhyRLtD9IJAEiKH2zq4qHNIw4n7wTl4Ux5mGPpv753hWnNbQO7hVHralT4ZozBgQxSjBo
wtZjNwdLTJ6kJuCrbeHuJxlgZKJ80dBjM/AmUQMNhzKbJBFSM3xJs100AMB3QgVF9dqHFG65D78J
n3Ogsk7c0gz30dMk1fj+m2Vt+yI+HMHnHv3ntgXMn4h+sRIADBeiLOZs84SD93HM4aHgyMLSRI7P
pgDYbkVul0zJz1iPlHF3flWNfIoT8Nggysx29I9ONa5FA/gGAfPIlh00NVJpFntylsWHoFDzuknr
rGdYt5Hm5kheASG502EWjdK53ElyS4FqpfsGnrK8SNHJmeIkfuwtLta3g01NRzdibI/Pzso79D9X
j0KFjcNizN63/MfrcuvbO2Ujn6p5bdeMVx3EOkSzCy7md/13abVH1u8hSnkVhoN7vmwagnetAM+h
ZODOeXk8QaX+qfb53q1CwCtXqhO3jcmx+AkGmg1rJaeQK5m6r4rNfWYxyPAZtXf5b5wtPpMCO4T7
t2BjyH/vWVelH94P//Pv7IUVy0voJyth1cmfPZAK2gCrujnXe8Zm6LqDnZKfUxt/4Y9fBaQJq3QY
VnxjkJbEEiYrXROcGWX/VJhHfRkY4l1qOOWIhFG8z2DwGP7ZDp5ejQjuSCPvFbs20R+EwzMLmoMy
IkRqiZFaznUIY+y6FzAp8ZHB6mLRNgkexNHRcUmce2krYegnkUPX9bN2xdajwIuZNupl6ttBH9K6
vdsygJGvjDEE/9/SlSy2l+VFZjoz8ON7e5T5G9R53eX57Vs18hAaDg/gPp7HuvoQj04QHfCXBe9U
hRtoCynaPdK2QlSSx+pHjT42sOrqRujzOdyz33LyfwEwzqcLNYgyx6cbjV3lDgnTKpKXUxLlJlqY
POmYa+lCqaqkGVSQU/oPxyUI84xNtTKiwTOyBanpnvJXM+Ou11VVmIrckqa4DFZL6OLT55F90ba4
hW5ZtGIdW/uEFhQbHASMxoczx2x1kZVm4mzxFj8NpnKJFUivKmt3kEMKr3foG0DV38Si8q3s3YDk
ZLdALcudFjxT8TsqmHni3FvzvBIlvWJ9EoeBWVSsOd4NNcDXq01tI68amQT1VlS6Qf8kMKIH99jO
9avNo/II7K5PBZz8shCJDkkf1CdEcnrqemyvGlmY1gaSxXzOtJ+O45qpBwQ/Le+ts6huTTKMIbsE
AJpDXja6aVOQkYkUcDM/5w2L4r9wrzQJXl3Ynz566R0o5hVLEyeTgEG1VJPErNv/3AdEqKGQ7w9p
QGt0lzXze85DY4j0+8vFnY1qh5HzdJ7KhCHFOQlvHlOz3tkNPWVFNqlMQwzioYwZ1tYqONporibR
6gVlHSPhON1GYxKLYlZ7gSKXqjhiaB8Jex8GyCx0eEQYcwDi7II+pjB+dW1FacuPpKQ1h+3B4FmM
pxKOcVk1V2UazLkLUT1k8STXvrvvoFpjzgjEnQtSRs2ApnxuhIpVgH/gMnjce9pL+E+ptH9R7nhB
X/03YW0o1ozPwfd/18F22zI2zTWW0Xbjy8qFGUEidYz2qfPAZuKatCmxP7qZ6n7AQM29jo+WdaHO
H5yXOlG3d6kh/tu4nsSH8xE0fi+QEQMVhSQK5mLKe7TrN81gu+OFFssqM6RY5CXTaOI68MbrJOdk
hHA7mCDQCn2wcEfezbXXLoQJ4efHx56LA4igEVpUBBYddjnkpato4x/zinsSH+Edx79REKBudnTL
cKiQRvYaS3ScFmaOqm21E8Fhq7L1yLQV5jR2YRTytLKjh/rRKKSDGuL322+0+kxMuarVPCZcez1D
U4pEbILzxeCYY49aUypuRHmfyy9dv5MemJS2GUZM2QMy9VPT+undERBqUQ/HWZ6omiQEozh0dzvk
ENmcoYfCk+ZFzcOc+jcwD6w2SA+wJRug8bzxaE/rb7E6RFVQArd89gUhEozqRBz/7v9OuZK2MXPg
izhiwnj2AGQqq7TooBJVijmaHsLFDyCfJO+s328tq+piDqHrIsoI3gI52VPybZZco38aWHBLCu5+
K8ztiq5RVbWhLY0eI6YixiSBM7eHQzbUDS3qOpBNvsqiJiwdYeuNqZGPdLwWRlH0UY0HOxXIuh/z
WyA6jGIahX3IGvIlhb5dqMfTnqNFGlBtrVn50b1P+KJCrT6VDmcKLUgt2YKKwvp8DRhsx8mHt5I6
viDYoqV64T9d+IS1yM03QVa/ASRIvwOWrxQx5PL7LH0oygjEd78rrrDaTrAjwbmyWWAO3G4meSfN
luHAgxxAwJ/5Q5xQPT7SC9un4qdz5D8eBlIhiYeuHYQQb2JLmMTreZqkgpBXBwBFRoKlN0VRlEPx
ZeBfW8CfKo3w6Fdx0sfIuJSaj1C5zsCLi+tQfbrWutyTy5GmD1KurySdYf+/ITwogVOtBve6tQCg
tfuC382GleMDERAgnKF0r13Ah+YK4uOcExgKzDp8R0j5QtaHcj+Hc8NB4Um4W1MJo10M0w1LV5SY
xUB/6BFwB2FW4e6ftk+yI+nCp1MBHvF8RXNDs2N0cw4yv8YzUswDGEPTy7LvGnQGkRYBO+ik8GxV
Ti/vK34ZPz19d0d3ZpW4PG29ElDdV7lDMhlg9Z/7B7ehUNhdWcJVikUKYidO5l7Eq+d0dFszMX1A
y+mVFNE1qIUZjNUpsnUdbN6Hr80YuMByU6AtugAChpDjAuLjS0BKZwSTOGV3WVAocY10btSeS/x7
/r1D2kO4JD0SzAx8hJNwXCentd29MGnQ6RZWd/Hudh82O8r6wiryQoFNzu0MdgaA6M9Wmk/PvWbW
WwW2iVpEa8hxKFKCMXRR3nKu4/Mmzjl1zWb7oPeEqFv5dDe6FGhIM021YcPPwi61WN5AAUxO5AXA
LPtK1Pt5wFC1fLyBdSju3ZgB41pNFUdbX0/AsbHjP7LvIFHh/qBDWHsSUWQtQfaLrAk1qvI3qtBA
n13EKkviVr7mE23icGsfkGafYHWfIXbpEv/nmmAnbdQS15uKs0JB3YOrvravQpvKjv/KEsh61X+L
6OCHtbnuqky7nc6u/c0B9O13XI6DL2Quls5Gyyf7GEr1VzJ4Dwau0U7t/kdE2xHiOhXN4XQ6AB+S
3NuCfpTlUhsETsu4UAHVDLQw1kDaFPe9T848u3PE9wzju1VNKFdwvbhMaWpYr7HL41rMaHlbuq/6
45wdzuFT9psddlmg6cNBZ7ZhWuv7/ULeLtHIvskAYHRV54PFMI0ABDWTXOfYRE+yBiv+CCFs7cQE
TIQPrhDZIRsLBDOcAIggYRhB1ewCJyo6yc/dkYNtw45wJDT3STPcfY8gRkbv3lIZ5J2fLRvk+XsV
z4pna4zBC76I7gzEmnHOyLBpQB8Ep7+sYQTgDhJqIieRQ0UCgEqMdXYDUzLCzbvJBQeCb9ltk5p0
IVBk4kss1Gv7xd6PQyaIk5kEVcNF0Gv7Wvlgvn4pJ0OzDSWd3qjtHHdVDEPC7W0w0R2fMkHgeiw5
DQMVVCoKZaYeymw2M07FQ3vAC5rq+dbkkA3RFw4tShg67cze0uTDrkiH/aIpg6Ges3QFJ6/NHzzl
xlcFPhzAKsy79/keaz6UyJ4zAx9gkDCi4/dCcy4NITTzhbiQN0haxidVEy0k6GiJ81YiWTqJYm79
X8tpnOdnO23LJKQeUyardwXve0lgnc02/iREFobwoNzIsgBx/1eHNkrtE1YX7AW4iUdlzddEw6ic
NDelk7v5ThcBMx6OHwcwjajc1DE8H3hdi5gTzicaNcktJm5nqijQqvHeueJ2yY0ePhxGVZlYXZ3G
tMtN8inOSlZ8t96CI8JXRQk4Cjfp0bqcSecrMeHJKZmXNXs64AJmrB6lFlLePfosq70Onqbg1dmk
O6aI4M0EGkjGuBacjmOZHj+QZzdmr2CUef4bArRX8nfA8HnefeDaYOY6+z///RS4ouNjoNf/JN3K
brPVuoFZ2nPk0tdEAGf4iele4MlZ0q5eSfwqZu7sgPssNal5jpVeDWfbDJ8TvExUQm9/YShJiSyS
RL6abyAsGYUgNHKfqWNz1NX1KCApEHBW3SWa7NkHt7eb+d/25rFbG5BFqIdPTS+dHjeTawpXitgo
CNdLat9eva+bOdODtYMGb1wwXNN5uwGEsOqi6sBKaJfbdX4JX69ch05j4l4JDquGfOFUl+km9diK
iptBkFl0jWSqRAaEjH2qSQHcuIbzUBGej8nUskSU1hb1gVimhDAklv/yYJAMkBv/7MQla3CLDaFs
Avko5TwJ4HBLjECB1E9elJvFReee7NY3brOc0XAgzNn60WI8wQ+SwEgSbRjttTFdb1+wNFblzRTi
Agn/ATanXDQ4YV4WnLMwss7/KCrACs18yz2GEJu+9VVNLbVo2AWZdfYBfCtoa8/oa1QfoZPKV/RO
7Zo62SxXrNdqqEd761+ja6c6A2+dEPg/GFpU1MYAyGbm5AWw/+/a6k63aLG8+gnFBR996Rdsylhq
rD1VriIE2lG7iK69ObbcksnRSDWkdzHhfTg2M4rzHWh+CwFx3jdYAhww/9B61JSo5ZD/H+DDu6oB
BfI2y9e9oxEJtGVG5AO/Ku0HjUeJU/yzwwdspRq05spDjCuae/LT9e7HcSnsBKKebIy75FVMlRaF
J/j5NX+5ST5m8mVldpVciTVPniZE8CsU9h6TYEdqpVtrIlJsGWdLVE4xeW4imo9FNmS5+MRqXkXY
EbshMN8HvdqZmMct8kTd5Ih+Hbmjj3gIx6BKP8BAmiYSBK85n6UFTj13MmY+rUgssU/d6cW/ErtD
v2gx2fjYF37/GD6mdjYAXDwsPHBfQW/SMCCoZehTk+9f808y/4Fdheg/XwznwoBFYb643NXpmekz
T5HVwGgJLEzJjb+GtiurmPTMSuwN4c5Gh91s9Z01Uym0WsJ1pcelsv0ePCF/tqCQG9DMjKa7Umln
fxyj/bWkO/0yi6kFxpaqkAJMOy2uHtx7LhlFIWvh9HPkdkkcRLHtBqv/DP+cBXcGRNLgK05Lcf7H
5/+qBkXWZ3abiuTuGy+LCV3xvs2Y0KIOFC/Fscju+cHqlaCEC5PTNbJe2GqKv2qWUnr6Ex2vUNkk
LN4h+JYKvbztFOs1DaDpXxGPOe7oP3g6FPc/nebgOnp/wvzve77EUeq/atLwRUB2jiUihAKo3diw
r0Wr5QgKGn87Qu53iGyz0o9DhLBC9q1P5ft9JPciesx75mWSqWrtaKWPzOMkhlfF1w5lQ3qYWW9s
Hr5SQrSsgI6tUokmyW8CwtM+9VJjlyISno2UxOqWxhicbGqy4YM9D1pmlPjtoSC8VUELPW7w5JBl
sOogGAFF7ePjDNG/yvp/DDsn/MrS5TojE9vhQvvfTR+YnXnbiDt/AUZQU212yyVc1bbbDRxz1k/l
V4/IeF/NcohpHyUDIzc7FlW3xfDA9CKzB9G0za3riOU53MwdX4bztgbR3pdf8PaAhvAbQjXbO3p1
2keSRN7eBJsmTmUzhnHQW76yPiTKEQq5lVuBtyV5YG+FZ9lgVLrS+ViqgmF0sSHoyRzs6WJpajzB
z748pBhXQtaMWtJIrmUxYTM8jxyXwtsWRz/kdOL9oF6LhAznTscfs2sboeCwxzRxu+9ta/I2sFYU
TZ7UcfcqaKkOEdBM08Jm/ttLeSoXkYCHtvLf2+i1bEBdyIeXEfIxfFyAV8fZOdxnP5mnE8JGN4RT
+dnKTyniVP5TGjabBOHk1YHWam5v6IB1QUaulrr8nRZaxdmCoLzNgW/+Ucl5hs1kN13TWww4+e1/
MaI7ZExeSTjaTUNfe3SIWsmabX4BkHBMMbgeg/Ng3HmzzUIPntnIJOqq88xuB/3VUJyhqlRTgBQp
Cm4sUq9Je5pC5Pg65Q+FkpglZsKlB9kn5DAMAcsnxWsX7U0HBCcEDwgwPHSNgbhvAEWAQZOIw99e
seReAP6/KzeAWMSEdZdwZwo5UtvsMl62kcAbCJzlyIhig5mojGjSmeQTsAKFXP+3mpUrCM1aHnzO
Ju1V/J0SLF+mD9UfUngYMKdqATmQrBKbugQ2NnduspVMUEi1ml4mzuJyFbQmLJs09MYSE6K2orgt
XFJ+rNE+xPja5w5C74XmiyAOousKkU0FajfStbzuKFO6TQTWTXx/0ieIktd5C53L1aS6ZtFDFGj3
KlHNfIUujR22E6lBenYlvt4E2tjEaWu6e+3Retet7lUtmStEmMAYoKR2nrzYciQQyZ130uF061go
yfuoVy8bX1ncsV7tbw6XBocWOFjn/NiOmi6cwqlGN1Kk99b208RZ+z63PPVMoQrHIjU6Ojc5jUdt
rzRzQjSqsRd27Onoo40fZkfQmsDCdkeoFYQkO48FUD+VmZA9DruqGKQozWRgsDibT5tlXEm2LGUr
SKGUCrkau8cVeA3mrplZnAyaNS5rrk/rj5bhCD5GMYtSPbnDoQFjpS3vNc8QdpX76FmGL9Qvv/D5
b/piuzMy2OOi0pb+I7tfDj3LmB3kkSjcYfxrrSGFb7OQVlgAFA+iV9OJoxVGOhftsVCgx0p5cKN7
b+bQxJMWPEOxq9cmRazCSnZ/Jf2pvUSw/ifWNQgRt4e6Q6DqUbVNuj1DibkpY5G2qVYELKJsv/4z
FDEnm7AbHHtRzoJX9fzkSAfXuQLyXLxiXPrFMur9SmFRG94f4JZVqkxbRrLAATzyVl5xtrwkUXmD
EgiFfv9U1lGMh4i2opO8bxeGj8R/+Sanc0gYOtnCTLp5W+xenrg1vXiyisf6tUBCYCZNIDCK5o60
Nk0aI0bi8i3UbGldjbsZxi7gxNBjxLknAVl8ROax5nTjECEtklHh1JK7goJyddc/BUWVJPtRY8D9
2iupK2jhyliqe7WIJZnq/5vIXgvJB0KwGJotlqACvqTR4bKvbXYxBbMHoAuaEINrdVrI1NVL8uAk
bbVKu2P3R0Ct/B7vpbUdlNAuTSnsPw0bX057qwXl1/ynxe0G3j+Si29sxJIx6tzl/ubsFtEzVjon
cHa6WfQZ0YAZpKOF4Bq3Et1fUAyc0Y0CO2aGOKtE0vORUxv6ohuJ+5pjt2k2zE69dEf/rn7PcWdi
D0Qqt3Hy9NnPSM616Y85xkE8BSMhflpBdqGgnzEOywPi74IJ/SFKs9IzD5w3aJ38DD7tyfqWqIw1
etsIwrr2+HDixf0Y1kUmvHznKOjz+26zBUPPglkXQLtZW2Xofv1LrgHLib+yUjKTGWk1pZvXpxey
EfFzOOtCMI2iRxXkzmGsKnzU4kFcJtF7yOAhR9TUy6OiL3lgUBT6ZYloABHewfaOBDEYVLjOVFK2
wmawy7E/d9pLwKoLCIlCq0s9HScEAZQWwsE1BHjSFaDjAllgw6k3dBnMl1e3iUi4qj6pDR2AO1q9
1tlUYkeAdQvi3z1gX4JzZpKpLK/Gjr/a2zNV7YW4/zakStePy5bw9Bhm7zufWMGWYfe7kHMqVMJv
snODgmauMs5PvUjIOAmdmVqXfVU2zfICOCQlmVSM+XY3QYcHn65wknWM/+0aIEgzb5qfGg4hwu00
itM0amP/olXFmixzPggov6iwH0tbmpWHPNrpVKXsHW0X4yIBXZCyHcHcEVjx7wXy0UVjNE9MlkHr
3Sb4FZTMZr+uMkD0+8EySQbTEqDkgkz3uRrpvWGBLclLQrNDPY5vJYVyc3lIG5bjo5/0O53hhGeE
o1kzK6qD8B33dP0ELa0dIwHAPmdTgt4uIa3chwaTaE+vaDYyO+QC0QCXdlCcVpVcGbIXoF8PEoU9
qPuBwJh0Bhs4MDZB6cgTBAy8DpfQtA1wqmMzw5gAOcjaq4iHeTWFKRE17aJmiX4S3+n6/NPmlJv/
Lu81fJ0nQ4bhVjmdW0rime8q9zLMk7zeHZVtxonxgsPi4LrHVcdGvAGIveYLqiWwwBvQifQac6s+
WsqFUSVS4Dk1kwmtTmxD0UdymqqXZazpLLtIc2sFHAROKaLcFL7BHUkyHLKRLkW9t/pK5bqBRtXh
PxSG5DE7yAfTkrp778IboiSU6pBkGUCDbEmN9ZQC4fn0VqRBau62r8Od10U9HM7IvCwom6tLbKdE
VE6kcopFNe0dGlEvfdtc8Fxmsul9Sp7tn+5SeTCG4KrYFWaY7L4rH7SGzWYw6RFBtTa4GeNMGmZd
PZ4HPvK0wRkD3YJxP0s0gqv2qyx4A6HmLSjNFNTk59ZgsBu5ub0sz5K6O9V8UEsSIMV10m7JPE+S
UmWUoH0rWLPOsKhYKw0b80eWmZIOaCGzcDP5SWTZVy9rFK1RwntJsPROJLQrOrWy/4PQQ9oDyHZo
UQz4zMc9PhnnB3LLtU0+QsqXOPrt9E0IGZl4+Qc/Zon/485qQBP16pCU0KpeQSkfeMorfPM0cmlk
kgafPXmPl9MIy+v/uh29nu4ZRciT4tFjsoHf5yjFZ2engM2N8Rqr+rnGKX4cKkl6U64bb9j/LBkK
7UC/wRNFN9FDMT07EPR6OMenP5Rq5oOYQyxCWxL6cYYpCgyNMF7Ify4SJtjK/agR3fbJxbWbGOnp
H+YGjdnjMX+MXad6mWgBRoyQLsQyzH9gKRt9L0sGCv3oikGIlfDhtAgQ7jcyW5kdZDSIFts4QDSu
vcRzEo15qzTTAOYlW0t5ubq/3TxEwixZIAOIb+zWVHdg4Y7iBLzIJsGSTsJAJUfNY3BQFkb2yR2i
wgBG+DlPNAazu+eyF6x2G58QPsvWMfj8ogLxhhj3mUZF+J21QobWFCILAScp5kkbCyKaAjQEh3/g
6+rXIvArhoi60mz2/dO2aMFNZW14jv8EoM1Do1Xqbz5urwE/es3JLtlWhQg4W4r9jkgjXThOGRzL
63b+pVRhNh4duqxk8N13tQFgYEV4lyR1YPJ76OTD1LwYa38KRhjc9/LvAatPBL8ETVrOjTfI6+Rr
Odrr9TmsLmq77aAPa4EqAUWw+jxF5VMskAOXbKsHOeHUZYZAoIodrN/NVzjkMUC+7E0hvFFSkQ/5
oAhWDd/ekQowTTRVHAfOsaJVO2rnBaSOh9QWMQSIqhxtf4b4SOXFDd5HT3FzjTgB5jHUIhfsX5YK
bwJHacbtMmzGUmpupkrt/eEtyQJO6w7Rjg/MFoWqv9QIbZx25409u3P5O3Nbp3HWxfaA5RP4qk1v
2ubL8T4o5abckEHTRCaUwMDypr5tk2O8fmgBNojTe4SH/PlyikYayrFWqGYCdNfSE6JiuYlHcwAn
rS/0a8TAM8BtYhek+IoEj944obto4a4lfkcCn7fm5s66TgRrBifl7s15cLKifr4QmT2psc8ULxFq
hkE2IFex5H8YMi/J7PJpTDraJY75Z/4fYFdFyQDM7raXqwWUjHlkenUm7tv9GfnnjmNDxR/r8f+h
0gZJA1rqVnS0Z/YnoXkVor6LozbFX4LFHN8IylNZ5Qu5S8IanV2Ay1O8AVWHMe89yJYVWhb7CwO9
EF36GvAtIfiUwfJtfNP3VgBes8Ps4FnlMX0dOaFLidiBr/2XeuVaf9iIjx+8e01slC3f+ZJr3MMN
e4mi9VWBHN3V8Yk9uVWY9swnvCrmzWOJ/5nmta3vynpC8T8vIhaR3svhrzZTGGJaIPh/NMzbsD78
zGvXxWSEgbVehdNIElke6H+Jqm1ElwWIxnHLiNq/lWnD2Fw6BnsxTTLRk0Qw3W9dIhvCoCAm2MjW
AhgYyvbegtIsC43YPuxAZRbsnKRy
`protect end_protected
