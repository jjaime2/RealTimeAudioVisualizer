-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wBLdh5nUwq0gNAAwJ4at3Z7JFM38TQU7VC2JvUBoUaFZ32X0hbV5YMnBdF+Xgg58Zd0DjfL4Aoeb
jJFBgKyo9eCV6IEktvnfMzSjVghjbnIknTfF2tLDzmvgnq20DuwNTFZOVZSw94x1LrzUO5BcYwz0
CY2pVAJiGXRmFbVHFKlj6a4ouwXerETHPgqZJ7cUJahJi9HB+e02ns/K4PtpYRpfgZ6FI0y2c9p4
801f27+fWj/87yEYcGQhKRMs4mghoGVcQufjO5nBCdkc1/cnVnTWyL/JC9xTB/OezKlGXqALiQv1
zT2f76Ecpy1QHGzzuUsLg7vY5cx0jdoCJ/1vnA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9104)
`protect data_block
fWBTXudsaJZw/x1Ft3zp6cxI0/ydz6ZbDTUxEW86NRJ47CmOW4/QxKMfOAIeQ4HeNCqHgM3XGEiW
AR/qfnhwTCDBWR31vf0ypaGwHHw2uo6dsNjjvFRhJkW624z4jc7/4hut4Gn+rF24cSm29KwyH4mC
nin5TU+gh8mpRzV+LevKva9R3LVyEYUkGBX1QYmC6YcwmEtSFWokX0Xut29ZIDm59l/SKfCyutb2
VBjO7lOtdUfmQ2Q8yNY57L4hMFN7Ao2P68C964EjGU9n2lnUaByJNbqOfQHrqlYdXoytO3e86Jc4
FFXzEnSsqAkIcqHQaW/X8nzIaV1DRNPZZjDp4Sgv3Vg3f60Al0ZUmn1nBH11m8Mp8vsatBdXfCD+
eYzr28gdYCtZ+5/drBJWilF4lwvu53Jalok242esoRctFgsqm6QEvrCOjom9zpVhYvedIThRKWFj
+qb/qVBobZZjUCk639ECeNk3SOKdQUwwqyA2d7b9MMQK/pd2o+93DK38FPMnMjFIVvzQbX6aFobu
9U2Fibs+ra5VVpCL57B3zgVBe7DRB9lZUobpJdraQXabvlEcn2CZmQc9txZK2plECX0z0VdSfgYA
uSKppVOKvbUFxQWr/6aVFfJU6XvFb2flCPpn2Hxz9khaN/e9h7BhsjshaWawPcCX0UnTt8VokcIN
WVu4MPK5jmKiZ3UAdY2lwP7VREURmgK4TBC4LGHzPZeuv9Y2xhg9+4nefcG9jsfkZKqYkuSXayIq
J3r8AW6XBecsOFjTBIo43G+G+MkciysHTYXpPGD3e0w1yfHVv8kPte9jl0ymCglrg5IIa2tOMwLo
3TVqC2PomcDg3d6tFiPGzHZAbTovfXw6ht+j+Ywtjx5936bKDox/iTA6o91v2aXiPUk5Ep9cn/kM
dUIqlyMWV2qvp/JD7NduVZf68+16F/mfxxEch9BvcV3toUjY6RnYaNYA7e9eMhTcGz2bwQj845db
uU9vgNn271iqdF6bCPL0v6JeCNiVBStSQJ6HDeS2nQVnrvCaSGQ/6RLkscx2gSrzKVSGaADXsldO
Rsjk2TiranTRXjn98MgVgGrkfPDYauRiVsYIV4WMIPdtBrmLTfeM89jlBaX+Fyj1ExoAODxZBfMI
t4464Fvq87Ygtb1frQ7uNWZrpTahNiLgFrLr3ZLh2GCaUJnkSzSCb1oiQkZbgJ23qmorz7zMw41L
7uIxorDs0rWxbceDgbYIJc99oTtCs+pjcwlilrgFfWDEr96FCvh2m4+Tz+F/GuMLGQFAqpdBG8D0
DF79OGZJIvHsaGzo6JasK9GfFDG5tdS4Im3SNDRqsoH2QZNCNguRoo9VcI5hKER1U+yeqviyK2wG
SEUXZ853JbkiR2/1a/U2lJyAGofLog3GrBqYtbsKS+S/CjJt9ND7HfzY6RRYdVzz5UYYyr5e3Rf6
EorNygq9upC8KhvZ3+vlFQR+4fmpD8+0AcpVqcK2vnSLwKqB6iPnwZ65mp+tZO8LY84T3X8C0uc8
KTzB2OxD5GimxfT6L6B8XvxO/Delnk2tPzJhh0xuXljlDMd+mItj3SFKgbFKukSwrJmkpR7rTEY+
u/EPMWyPYewoBgcRnVVbf5vzDce6rLeGWipQ8gU//kruxIryVJANu7d/H6x30OBJFuTj8RDiptCq
E5ZMKfKRRPzQLo2rPzxUWDbXqIU9stinACnyRWfvNfh3sBk0XDruwMUhkvZd2EXiWhtSkbs5sEXK
tpscSReZCD4BWLju5Ub7uGbAYP7twaHeu5hYSHoIWxoi1Ujd77NN47r2V1/rD1jUksEGU2asDZQl
lIqbzSU50jvX2mzKw8zNvnsSBuh0vnIe+BxACcHPBd7eCLNu6eZNZqPhPpPoASUIx10YGQ2UYu5b
W9LG10t4/g3t7dW4dcwUwEgMzZDNLh4Vt5g8zP+YRiD0up9CuSFfmXcu+2d/AWl9nLmZ9yN8DN2w
rwZxkoE1fIbgjTUjMDV3lN2Q63GxTZtipcnewfRA3dynpz7OBqRgfF4GiQGl5MrLd4tDaq2TilaO
2XENrQ4gmq9Q7sb21xeQFUXNnk+TP/iepSsTyoAMhQwRjT2+uLlmnrrOtklAmXzv8Z8A2o1pl0To
2oz+kmO68+iyr8skg9TUY8ECBN/rF4I+xIXLlryuyO4IJl9fiIBl8PpiwMiANesz5Q2lZ90XZ6uC
DxgFcEXLxBNY74AK4V0355YlnQPij+dAA/btjSnx0miMG53VSWd3WehvbK8jqtt7+khtRpRP6aga
GFYD8eCq31t2+qF340Lxo8ygtEcFR89SHyz9qlylg0ABhQ1JNJotom0Ed7m4Z90T6//foK6Zfx9v
PwReMOtBtHQswhaZVEzz16UtUS5EhBipL9z1OLYLSQgpMqoynzEIjgINmzSlJLOHWhs4g/njx01V
yHNOuxO6uxSEXylUTbvsAtpsfI6i3LRCUwuU0crHS6+yjeoo+cJub/s0tc5syAB2E06nwDIvebL4
8AQBLzRScMtGD+a7CQN0tihlFjBUvnUCZfrnL8g6GhDUfudEm936+UlWbN9Kz3rGTQD8DMoVBVVo
KBZS1SzRc+vLxgOry9ECW2KM331FHXAcYZKjZFui5LTMs0TDzDyj7hjmVVdfgDyz2Qg4meht1Kz2
zqnX6Ri9MdWqrnsVvFCPJvIb1wQ0kIS02dev9CoNrc6EvRtYRk3WLpdJm44lSKszvl8ZtViSuFD1
fy+G1v9KWxUG1S59U09g9KCe0qinlSRXHAjPLTOUeJvQhSTzNfDvGnQBDGxG4rxMmSMPE8dSbig8
GcKbRPD3nMUBNqjATacTZpuCz2yA8ob40gk283jgAOfkXdE+7DHPALdapgtEswDL7qHf/GROV5F+
hNMgIBs6P/gB6eY4GKCVhgu5U732dpNEK1xa6bBc160ZWL7QFwKHF2ya41HKUfSOBFGH4HQ6BWiG
1RRPKkohhZwsjL6c5KQYjYhUMozXEqxTcZk0UnapBI+uplbSynNhfkb8KNzjGFGK+6hFZZk8+lXJ
q4KS/MxTARkPpVMXgPYMvOZ39zFg5njoLLq2hKcVj2sKNGQxb/fYs0arzqtbEb17g8lBJPRY09TD
9+PrSoOTtBr2YwG/WpPdDSsvtkoibLJmBG7n1vXil1Z0peJhONs+P+5pkt4nJhXqG5fMyMtkzsyS
Fzq4SR9y45tcOFaaHP+ahF0n7k5P5fX+Z2X/rE5clZ4KbfEMGomAK1Q4wQ+/u5ct/L2EcPURvwSI
miTdS4t/7XjzaHm8W6BQETt1ZZ7xXXh2SDgrpWV5GKaV7CjpLiYSGTGmb0S4DuS3ek3MJzEsh2vb
4vVvR/B/k046I1K0XgLn6JpxijHR11Sa+QbDluK8oxO8C0jmUjsJQyLw/cIN9ERlLRUt166D0r7/
Ctn6myy8aCLQEPkvB1TBRoSzDEzBjSAgvfWFeAPAF7okFfdKLdDuweTBTL4vc3O+C9kFCWYtZn0S
q28anV4ed4F+RdmnEfeRCPIoUiD+khko6lgC+FaHSu3/0oPmiN2sRL9zWJ1LyCdXM9Q6osZmCujN
S1YjfkqfLbOpN/4IE5o1wn3uuAeCbYGgxlNIXPX/8yIXCEvLFoCd2fx590+e0Q0exYCb7mfDoTyT
oo8tU8dulEVRWQH1Hr2SYp5VqFNUj3E+1DNu2ozOACN77vDZM8ef3w8E15WzwtLIOJ734Vwon+Re
gQHua9GWHC0og8jqSFfqph0YLIf4PWUGFsRAniVG02RJQCXqvQ5oTS1TfDOCQXe2ez7WRLAlFmX9
0662w0BMOZm1PzDdEwBUGFtavrev5f/ldmjUN/ux9A1ukKXYS+hR0G2k1SBV69/xWyIS36g3a8nc
saHqC5I3L66oQ0V2WdbeMYAsj7qYUrGYzBWGrDm38jKE6cW/8u9CQq35omQ0XsSCQYBZ/H8X6X8B
bzITU7k8KfurXrGhK/ulRSdCMV6Cw/pmUr+3aYRL8+gH1u29Zk7AAHVU4tH1MmsbGVZymfekFzoj
a3gc6/pb78frwipQv5MhQlDDHqzC9RZxhNWqnjFmT04CZqho5mC9hWzEDOteDW4hP68HnU6ynF2w
b3jQlKxQ72nesltejQOCy87OUlmWr44yOD7jHVrtgGIg42AfjyzIlR1x0o3v1+zm++f0tlwIl5I+
M6IThgYj7yED3aSdyinj/T2t2JVWOALePm1gQUwX/I7VjHvxjdlLolIRLKQUGZZjLOaIe/UVx5lT
D8WO9d/AbU9zcp+VhPVc/0Rs/koNIHkMhPsGOOiiImhOv7Z6N3b4GqERg3cpXi26FeIr+vrM55Tm
DhpVEZaHwTmo3IUggXTcwFNdXZ7UZXFHnAwB/VmFztpHLNcbOIknd16vobj7bI2BgYKJsmYqBTb+
FCc4f7JTdIYTvKN3aoN0MIh/aJzOaebYTN+Px5HH1IFjLbWo5n1QbxP3Wamf4bF1Qsre4EvnsYoS
LQbJx0ccnzytuwULHyyYSu7VQJOX5tf8u9hFdpwvWBaMLrEYoydHGg60AZJ6j7TcfR/QzzxJl4li
YY7Q+NLQESjxBeU5Ce4MT5q3FToumMRISyA4aYPboWKuDzc35b3JoL7g2MEFI95lW2VT4V7LHAlD
I7XDgLKIGsXBz1BbGIY44K9LL8p3Vt/HoqOruGgWiQjJBGWUzQpzCl6Hi1EW9yVsz/yfZwpq3ghu
MnNntPPS8jPepRciZObjj0hrfNefiX/NvwUjJSjYK8zte664gdKHRcjWpKQzkGKvNA6BanfoAsg3
GjVJKAJ4l/ha/o+LbAcE7tYN4y4kF58QSArs0XMDP+DCEprxmxHJZ/qoZVWSyP2aGN+k2CyVHZg4
ZRRMpwmO0/6JOC94qey2UUpGcWD4jaEPiaKcYWq9MpNoOUxhjdpN3hrIsP53hVNepWzZbFnE0Zw2
GIevtz0L+qivOpay3Zh/QaKvPmVIt3fDJEkkLkgk7XOKG0RZ9IUjZ1p7AYE2dnMG77WVmN1JNJvE
qIBimsbOoMSDw6pJu9mAl3e612B0H903Jtoc5mErsKwFH0/DGInzUdTK6mvYF8uW9o/rgnHjbbIC
Bs8hhZp/tCAHQG//kqq51N9mAuONgpU3IalqGN+9ofayj5D/AOX4Od/G7Hu90U4a1FGueABcHkt/
frW+0l1Soqe2WfWPx4B293ftkrzbAja2JJ/wyt9QX8786jjPoVPF11/ETvAdJ3KZcR7bKNWrM1Nz
+PSLqNvT59yjrVk8yovEUu5HKeeQIKXrkAPvljzMMrEUlLc3LEbPB8xT+O0alQ63BpaPzZ1/bxL8
SytY+KZzyy9clLrbVedZm0GY09SgVNIid5CBK0hULEEsZwf+PTvjbAiTQUNQ6Bnyeo8Cs2WWE391
whaEUgZF/oSXIGs/npva8cQ89ofa0UuB2YNtXUULPjgHftfZwm20ijZvIAaGh06r30C31krdB01/
/sIMctp/EZbxN5DE5ZGKsG+3eimlbQC10xFC0W3k28SX+lBZ735D54TQQU6KRyChYSMxuJg8qlHH
KsgwF/McSyzmAWvcLY0PKgancZD1FTwANuY0hpJGyyBa+IxvolT1F28IVmETkgBh/PQ32Sd5WH+S
o4yarnjnWHbZk89XI7b7jpU9sa3C14bz2beYy/JE/Gh1jesl8dQr5LhiEm3unXog361Nat1NL15k
ZGsbY5LHGFUmocp604QHCVSQ+n2GDOoI4PubrkxIa2PR7wYo6ArxtiYlZFcBZttYFPN6kN+brluk
lxxXIa8C82ETuRWDLu1UC4DNOidnxtvQR56D1tFfGCm90MwqKM4IPtWSkZYXZP4C34Hk8s+svdlu
KC8K974dZ/5DD9IJVI+MVNFiacBqy7j33jKEpPqjKpVoy319t6SQTDZ8dYmo+k/PDgIczVa2t5vU
sNAGu40Y9/5noaz25ehyOhPl2xjPFU4imZo4Uv16rO357IGLcbnEJoEyNEATlO9ZZXwzIjF2pYLj
xBbPrW1Twtw/dbEH/gZxkqzTP5IXSI8CuIg/iWRuWxwleGmms15YWwvdKTAdPXPh7xrKAdz9KR37
mvfTabbxR15dhO56w8HZiyKeIFOKgdCUZTrPLvmjBuArXAbOt/Ng5tfkxJXjkDwA9m92TBn7mINA
LhktWhr4hmFAAF9r9UguzT9Q0rxZ3fLLBaN1/lSM5B5mSHsnJE/eAGdanehGVcbRTEIW+rQLFxlg
NlRo92fVmrIpj0zPYlwh/5gwmEoXumMq63cvGKHHRMv8fU1Hvb+gOW+JMxmOkf2c9ZDCIIaQ1/1X
D/H05w4kMR8o0b0b1SzPjCw1TAA2daiNTm02tu6cK98PVl5rnfJL7Z0s7PHMG/M7N6hw7wPPpZIB
X2CSzd1dO9wyxl71ZJIjJgvxsIY/ighHLJpwnOtPWiYyG9GhC3LYObEREQ7Es2mLFE5THJmCtkvg
Pac045RHnI7Pkuxfs/OrRRUOGcpTYy1/msjswicuvtWQpOCDOIuMKrbqEVBo8zYPtRDiti5ajDNv
4Ei4l27yYpYNw7bpPoAmTwhODAZsX+knA4gDJIoUoyBtTcI5lLr7SRRDBlLCmNEZQ24tIChFVYGr
8dE6/CMn2hFDxnZlXS1WZ5PE/vrS44/CgG8jD3EBQQUBKb9FXA2Pa8oHVjGLUtt+ZaziUYMXBbFU
EW7DCVHWqM/iV7WLThM1uIAn5IWqyKMDSY8F9CyyPbHGVNYThOfaIbR99WrE2ibV+qV8tUPAFVtG
Ta3RyX0MW4w8rz2EwysKdVF2wmkAEuwAtuMQBvRB15MIDAynCq/PiRV615WwPKZ8F4bzPIo3GDbe
PuYgs7i49XlHiir0l2l9l+4jOImbmPO1pM/lo0xf8Il3blvTr3dOofvwOjr81lqJ0urf4svpq44S
QQlZdyHOpV/GOSZ75JUzpdiYLTI2bLwe7cxJT+Joaz+yD3Ei/MiKNVrYeffCLzvjQT+hkMHDQnLy
u1mPB956EjOFiZRR+zk4+Ngndt+4NJqdhix8piyFIeUh/fl3IbTj3zTyvxjsYrYtwK8UO9pG/r4m
mKCBJMzgZ0QBQqm1Y2bM0YsZJOQ8Kf9BYMAtCLpgeY2nuZdgM5weMP46nl9tEyBHutnN5nwsYkcp
2FFOtIiOGlEWGAhMh8QXJx0w/Z8OkCzcbHuoqx3L3CnXusn/DDpevuNnzZS6ufHGr5BZkcFSFOrg
BYGVDYRStTXkpXFRNjw1kskyUD/uMbDoiTFFYqmt+p6F5qpagXdksHUnaJdtsxFmBCQ+un4OsVti
FxlqWlOdeT85kJy1TMJNEa0Ub8RUZRurJm1q3C+642HORo10Al3aUX8O1QeIOGzp+qj+pGMxSAwk
U8bRQS0rapttakvEBYL19kB/1gaIIM9g+8ubxB3SQzFUwrGvgqt33jUgqWnpqnBy63RZ2LsbMwPt
ccMyAH54xx6MY69LXm0q9aEACVyNGDeUYZ9YfrLwIkCc0CB2dPRbBgT3Ij4PXjisA8jbdvkn91GY
bxvs/4jpn1jBfA4XcWHzI/7damQIRi9jNfc8Tpf0myZnK+p5fKF4GDpD3lwtzB0SCZW0u4RuKvBr
pOnQ+CtNfrlBhDVukd2OKVdu14l9DJI/7EZCFAb4Mo+HIr0gvqmayWZQ0pX3uen6jE4093QHCaiQ
vweD4Pdvhz6MwntyvPOPLe17cZ1ITWLP5f85MXpG6o2Sbw1LXCTv6Vn9fm+m7K/zU8UbsIb7K0x9
KNltNpp0rNa9iDRsSbkeMfaWK4ykHxKX/kR1HVcRPUrlicGdcYLguZBepZOa5gCsPvybH/s1nvFm
3u5ZLz/ZAIkY5unZ7xjqcmWiOyVZEp6wgCJO7QjGrF33FuOdva8xfYY9iKhceYdqdQQ4Kyd70V9v
bQ6WKLWmwFSzD19crifFYGQlnJbxHn5w0Ry4cZ/fS1bjumLi38+mrVjVlXHGZ40lqItH5XEAL3H6
7ARv9QaGTAPFsFDlO65qObdkwrFRCWgZ2dek/+UykyYADghBjdxqNM+bf58661aaTOycv481OcIV
wmmTDYoIyEdWXTlY2Tz0H+mhIixUQqF4ahOeJEMeDfIT2fB7arMrcpNtKDw9JDzSSBriLoL9hQpU
Ze02qPm1S9lHzkcEQbnC0G86PMXUghw34K4lb4dJWfkFShAsHyoNk348PhYvuk7QGXsHh9ze4yHT
EF7cBhzDV/o8q/kXZEaKd6YxH128aV6d+yatr3wz6Zvrzup9UiQi69WM1wAeq38OzeV5lv9IStgN
F7bAkfCVRbAP/7de6ndMI9vbT7qae53O3pz2jZl2+6CxIpIZS0rxls4BzKiixiv0oU2Pn9OS++aq
XdDNXn6yBWDfyCxc89rtP1xr4cBN0hB8NbjKaZgJ2eH++I9f5aCsFeFMvljBOiaCBL6qHr9j3WDb
x5NLB5Gy1sRoGi2c5H7TMmZh1W43jZsvrGItMfSZ5zZFQVaRNWlTU0GcHTyjVEjZPY6p8/rOf6i1
wpdVAJWN6gQpJajWQUtUUQVcI93rgw7Y9GCjiAhvHZ+rjrX8JNLmcA3Bm5e5J+Qiar8AaRgs8wdz
Stx+YKkqvOn5sxny1v6jurhLt3uPC5GO68ZIkC6rczeVAgGVlwkf3dE70JOaZNWIx/zqd0exXui6
8V3a+62LaDiH5HJPe/SgvyaBSJZ1/WdWG1g9En8dETARfAOYpqSlxSnK4ES9ZiTbevEU0aNnzOBb
zYlYqnvY5obJfys4bc8UXeArpljCIv4Jww3FUlY/G7nMLK1dgKserh73koXkjtO/sw1zNvK47dJq
4mGY8rThhLE5RMpXTDWwUAb9ay6GnLSJr+4SNue+dz1pE7DrrRICa6zbO87yxmYx35wgosZ3qHsM
rO9ltmLqwTd/weJX1kgoGnTrOgELwTWnQDJc1Gmdlu3uF6t3wInCdj3TFQNR83kBo3JdZwg4d332
bxtlsNd7xgoTOKPRtwQ8pLQHd67m52QgSa7dDTMpo6kfuVJgrHeixJ+WmG3cuN+iNMqFWUQCtXup
3SALOWBxQ/cZb6NUY5DrPHaXFltmCdGDFgn3js5fCxBGoBeK0W1MB8U7b8Ld9/jPgvd35jOQXwOG
ju4jtBuCTFK++GrvvrVxwoC4kZ0X/dpb17wrzpWYPRK5IDDoIasDKUaHyO51Ds+zOuE0oQKvceo1
M6ATSHwom3FaEB95mZ5bbiN0n7nPJh/cnOjJPNS5gBL2LwG+HF9ZDUJhOldKWz/XC6eH3/rpo0vg
ulUQgnKJpx9sDefND9ls3baz6uI0Bc1rJ0MZnc9R0uxzZu320gugXeo/KVyQ+ub//HRM4GwisN6I
HRJz2giOh4DO1tLxrt4vh4Wnfx29t9pbCtCxIZjYtric3DgyMhsU/6bv2Tm4KQptuhxiZ68FsmQa
eNdyuQ/OHQyebHUhrPGmvUklng+PnS4sneopzuVVfx1aDXw8lEVGQSlOhTaGZFBJXZAM+YUDDYga
2Oz4ONZU3e7gd6L1bu4lTm2j+rRw9mf64VdFzECKEoseycAZuJzP50zpDerIPLXE5uvbFaIT/8XW
1o092mdu+ew473vgaoPk29MqdWb29gVJVYwZw7jYUogToI2vQKgnVAsvdf4gFTRJ2zV3xapy9ZgB
iNPUA3n/aVZSrLjJA0ouqBUpn55GmHFdEQri7Feh9trv8yxNUV0dcOUzrDOPeJ6E54KasyDPT8ga
Gnsoigetr17gUu6aHg96nmd5qtT7hxUFDnd35UryqKZBQSQQqU5tH0rd+5fExe4mbklyXVScuTmI
oIE2WVgH+FldQjXWRFoc1om6pqh0fYqJFybGbz+/4zkc2OWQcRQkDl/MT2bYP/GitW2JhOuodobt
4OOeg/iZhcwLTyQNyK2NbS+Qh49cALzlA8CE/Pfl3HOPPxVWzHIjMKzBhyvd1Wg064APkBq911TC
x1GSOL3WRqdlUEDx/PojbSky2baYHg0gPbE7v1f52gs4HjoB39MsvlYKVMLDPywqdiI4O5CHbU30
tF4tGSCaqr5VQzVFGzo/Tcpt88gsENFx8AHhojHJVvqMNrFVFrihgWdkF3evFfIF8UDSjnTiEqOG
/jFF8av8LSUsvPAyPefA/g2XJsi5IOxmYqfgamHxKpaOJF2bGXDFU2f8nJKG4pemrU5smvX3Mo1g
3pAbz1dNpPmTiB/dfzjrvmacWHRyeebZB6Hq0xhbjyCz398tW4apYrpjEwRu2yR3XaRutDn7Yih/
Rp4NDTuJy5+f87RzDujuALifZSlq9QTZxW44y/y7XsIFE7vItxCYD0YdKXwDcgaxYQ7nmakOwKlZ
Igm9HV7EJcPKklRGenxUyXW91Vjn1w1AA/aa6S99JgZ0LYRpMAwpNXAsoEyMfJYD6VDjNn0TD3a5
Ok9N+/5v/Iv+58l88d9taJBYUbrfJhZn0aY84o1LzBLSA9UqlKtGCzcfnpRpcbEu1veN2NwH2A66
wjVk+DtmX8C+nUJa66NPnqvKYI+RnCiS1SX3BfYemLySWsg7cymeT4VPL8d3OJaO/PhmCArkoDfk
QM7lA1lu5FeYzIAh6P5OQWA/1ZBY2Z6LHMfzvCPbWDenlCYinhcqo+Kmr6ZfZuxJgd4g6MgQVyNJ
0WWPi7K4+fVGGoej9/bA2HtHd2MopvVA522+6tL8XdEyhoE2gfKP/bNX1V0TmIyZGRdoFU44jffB
xVVCmG0hXV4o6zSVwIbGvD9mVgJMbnSWHFHhrw6ZhJ591u5DFNYIa4lzo2e5iZ1u9FAxO8SVxUbB
uAWUYoFoPyYXZHh11yUawfO+GP5RzGIu4oBr2RuDBrXl9rxj/q1Ua0WCtdUI80rPOVpO9IDDR0Ur
4wCKXOAe6UKTc/B9AqUOAgK/v/fiWYZsdwOb524a4auJw3mb4QhDJWkKwsHSlGUSPsOJKB2Df7Ng
dGbOpkzIV4E7lCOnDCxLsQyNvKyitxTJYnIw+GFLU+Y4nMzmSU2zPeUS7sN7l8Tbi+CsfTZGUWCL
lkAiBsdKzmzJF8Je2KoDRgY35jeEBJtn0hI5mQ6Cus9YTwr0KmVUIT2x86opS8fhX3Mbnajlup+A
1c5P4K5AJ4QezcnobW42YF2Nm2uQRAT3Fk3Ob1RZe/ihFAf93H/DSDeoaNSSGi0TtTzxeu1zJ4f+
GtcuEHyy5zDVtFw20wVX1ZpFViNCbzz3ngyfiDJKmZh1xx9XzvJOoeDSZGaQPc46vUD7m06fPcqL
Q2WMOX5qSkz/olZIBp8jM02zJcAQE1AXwHDj1+Whf6m0sHhAaaF2MrTdoyEOaRpzTvKi8Fksdq5y
rhip5uvoJQKXsr6oSNCOVqJ9mccBD1Am5jtY1gUfYdUKvdk7ACQVx/yUhofasaSfkxioTFm2r+hN
CnnlqdtlkgrpIpEHxsbfhM+BPgr3cATrvbC62pDlmpMLk2COdcNw4ZeyFHzAwxEJWdT6bN3OO/Hn
RPPrG82YUhqiqh1css5N7aihtkmcYPJqNfXwxmFkIBqvUkcIn+sPLgR/IvK7aEX2Ene3cOsptatk
IZ6iHhUh2loznMJkNTK1KRFiAcpPcG8TDpUFPNhWVcGl5rUfLRqOPLAy02dbtLSe+3pS0SPDe1M6
cire9CvTOrh3wdhf7hoipHcD6wj9GvDj9wja8piIwCg42cDQ9Dc91ZXoDx3T8F8b6gIFK75pqBZ5
1CIFdoOsEknyHovgp154IE/AuVtzqe5TnByjBq92FGc1+xZZQGbw0uUSS9unHBV9wDYbRQefcihk
dLLP7rJjDepKrIv/qpHvcwhFCFlWMY+lC6W5r0ITFQ1buAIP6LOUEwKGci07qOWRKCYa225lG8w5
UiyoEixPjwfrZmn8xl4Foc0dbWLdtZeJABU3JDTWn8pKFrMSExn7blfMXSMf8O8cACl4Jh4bKxsB
9A+JAR65nFX7oxmPXzuvSzKKyEChcO1pmIriiNAfHFMDxAFlwcyNTwaCuH13+el5siMrceS2TKaI
r96Gpm/Iael5fVVCk/sqixq0a6UN2h+xPxmz/on93Y7wqTXlbN6wTbrLaHMuJrJ56890+xdRqAty
ikH/4MUkIxdNMsRD/qDDfJv7m5UdYNf2CyFFCA4z9rabFk9gzw+2y6A=
`protect end_protected
