��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E�ﻏ��Aގ�~ބq\�l�1�4QQB��t�
�_�㬃1Iw�$�=�\�:�}Օqգ�$�ZB�h��NS%`2#r�e��c��B��FJ�CH"!��G�D�}��_�W%�4����QWB���S��4*�+�P���Hʚ����a������.�CċW�,�ɕ3��v���^_,���G�k�;��Z�Kɪ|��5���T#]I���m6�{iuc� �y36��j��,�ٱ���؜9~����^����}��8@Mh���IR������%܅I��I:�/i\�?<e��!�gҩgkj� �{U�T���@H�K	o����0����D�G�D�}����6P�N��H����u: t��=��M>��)8Li�ȿ�g���mJY�7�\�}hsxI�@�R�_�=�C�xb��ʑN�| �\}ID$���8�gY?�<D�ۼ.{tVk���O.LUI��Z�`�0�f���w����p�@xA>�n)��0/�KP�����Oα��B���4雖\�.���5�l�=������9>���]�
�%���#C��8�X�-��>�.��ũn۔k�؁�QO��I����������zj�Q��*��ke�n��%	��<P\8�^G����4�c*��(l�<*,�o8��\�峷��1����X�!��Ʃ�q@L�<���np3����}a��F���c,hs�'N+;�"N)?ϕj/�y*�F��W�?�;�t�.�߫��`��}� �?��흹����"�&X�����΁�� j��㦎�W��~�w6UN���4����L7�b���l�sL����x6]�F�9�iTBU�!֚����}�=Zx�A�8��: S/Y���*1Č+�PiL��)SkW�Ő9��i��]y���X�
B�\��W�W$��O�"8GU���
h粒&Ö��a�kA�`��X�3�P��a��w�*kP~Q���N��}]~����AdÌ>p�������ɜ��,�Nq�l����sg�_[F̿���Y�����2�XA�A�[�4��mQl�ٌ��A��^��[ؼ�K�4j<D��+S'��B��0,����+D�h�p��qm:Z��O���Q`�������s�`x�j;{L���Yy(��Q����a]B.Xې�f>셌p�ŀ��3O%x���	���<~��W�<*�8�r�AH#�^S��u��)�ԁ�����O�:BȇN��V =B���
=�ɓ��u�Q�l^0sCb��C�m�?����$E��+�*?:z7��W�f7�'��é�ڣ~�2�4|�'�\�N��h66�6�u�1\~�����:Zn�Vx�2=B�-h�G'�Ơ�1oMQ"���x� �]�nGB��P�=?����b��Դ|�8�vm�!'S!�&B�=�>b��/typZ��_�Z�5���aI����+m;���}�I9�����Ci$]إ�����p�D��o���UAG;�86�`����F�g ��f���T�D���҄� ���N���? W�>߶�O��}i��$\����h��o���~�V��WH��=4@����|���I��s^U*i�XǬYY�obv��tXA�u1:w�Jv�'x��N~���)[(W��gw�SӲ�|�������O���be̮a]t�mO �K�>�~���4��cܯ�]�fżz�����YѮ`��t�ԯ���xYZ���
QDsr��M�3�a���a�%l"T�����G\ΰ9J2sxOS���)`��+���'	Y���Bh�k�moW��}���z��w<�7|#�d�'e���mԎ�.��%`�j��2�:FwPD�s̀K�V��
���#Eӣ�-h&����P��%=���ci~t'ߦ��k'=z��b:�2:6݀�T�jf��0_�7Pi�/9|i���=W���tayzA�G���	Ҫ�{��^�~�|�U��hH �6%��Xʛ՚�9�kNQ�4�-�<��Ǎ�+oyt��=߰~���7��~�"�3�BHW����Z��0Kϝ0��m޶����ɢn�ͫ^':����1�
�9��{ΰm^�k�[��'��nf�_�B҃�_�;��^u�=X�����<_�#�?q�k�� ��� ��q� ��P�H
�o�Z?ŧ0���B�J����53�ks^.t�M�/4�)�F6�,��t�yr�8��S� ��R���� ;�[Kا�����}��y~��>���C����%�^��Q�;�j;�_B����)'�Ws�oM����f�Ml��/��w١]��v�2�� �R��-�p�*9Y���3V@L���N��N-τV��pFh�tgj)�:�?�
R�J0�o	H��m��U{�Q�c�#�ew�%P��Nb�K��c��nh(�����*	�0�(���Mf:$B�
tj��>ת��47�u/f�[�=�XD��/�L�8���B���75��n?0ﭖ7��'�ev�˦�?�8��vF7����؈N-����#���i�O˄O�[Ƣ-%��Ջ���y#,vI��`,�d#�\�?�X �����]Kc�w��~Gy-Ľ9��c� q�ąO�1�����3�� �k�>�0��*���g�eJ��������+��-�A�G�Q�RS�`l�����6�f�?Sl|i1�n��3��2��+�98\���ݦ�����A�$ʢu����r%�һ�Rq�!��#�߉�5Q�,}G�@9���}��+n	85��o7��Z�I)#,�aO�W{��2,��陎�s�Q�ml�C���f3a�d��hXo��'��Xva)�azU8
���9�FL��Hi҈R����O�z��L.�}�A��h7
H�0j ��l�t
=��۶k��Λ�%�SB+��U���S����{~\�	�t�Mϟ�ny��Y��,w[�5p#�'^����Eѓ&���H�4c��	&Y�NʂŔ�w �|rP��N�Y����؄�J�-*7 �Ȑz��2�H�oe�����)�UJ�m��)�D��S��D�~��>s9@�q�n��o.�a�^�r�5��/,6 8u(ݮv�hW�'^��<�$����@ܞa.���zq�f���B��#1�d���n��G�D����)*�Fg�n3��׬ý�f4Jν��R�T��0�>�omf�l?�Meb�O>r//�_����B`�0�/
�8Q��T��Y�p�T�L���U�Yf��sF|���1%�\S���
�(a45��=tI�b�ei�e�z�H��A�~R uǻt�S@%�$�|��F�;y�0�Z%��݇IG���K�?M�);���!�Vpv�|���O0���ڑ�MmB�k���G�U�Є��?�x}��r�"a�hzEd�3�@��G��S�B�
Z��,�\8��T�J�;���)L_�c~rV/�<�>^�H!A�O����� �Z�zo�N������o�pq�䬓��gOtG�8�g���Q�M���e�,)Ɨ\D��)��"����R��"�)zU��{ז�e�ʁ����,@t;�3�(=B���g��z	;@�P�'ld[��0�KJ��d�yGd��!)��1��T1�k�"��1�!�T�g��#�2���]�FpQ}��@7��N�>���D�߽p�����_��F���g��Z��g �wN�KX�f<�2uZ��	��6�L��ﴕ�	ۤyn��`��M�sA�m����
-O��Jd1��;�����Q�ɕ_Kl�}���2��*¿���k�Guc�N%�3d�o����0���c*�-�m�#���=8�R�_�(���B��vƹms�C���8 ��a�p�W�у~ת+[:���N��$���vg+HS�c����w��7�Ԏ�=��˵�8J��e��ʉx��4W�t�Q2�����@ޏ�^8��%=��4mj��Z19\S ~�++�ƕ-X�2��0�`s|�Tg�ϕ�FVҎ@M������)&��D�p ������.�Q1��v7o�-;
���Ϡ����w�kE��㧩*!���$�Oxo���cq�?s�)�o�]�ٚx��R7��3'`�njԫ�󒞋�gt>��"�k����=�gf�0��r;���=p�" �fN�k��1���
W
9(dt��@�M4�qe�.O�4�ቢ��G��oXP��B�9�gQ]+�^��$��mHͶ.�1�d�&T��ޔ���%��o�}�F�Lt���ڌr�x���&�k�e�
BÆM+ܐ���ЩO��T%��ye £#K��.򣄻��q2�,{6�X^�A������v�jVA�oj�\�.�GAj⾧fo��O]�0h��1W��Z ���K�٦8��t��T�'�n;��~o�����&�D��$ʖO콲�"�M^��őg����$k�v�,�1��^݄���������L�Xk|/�[�dB���v��ZQ��R�R��k�YM��i!��Yԅ�	EG���A�*k�Js������;vM*�k��4_Bq$�u}��g²~`�t�� ~��\���J�vMPu�d����� �t."$�Q�B����}��m�G�w�L0����(K�&���������i���^�=�X���)=��2jl>���y�K;ʰ�V�Ԇv\�{�2]�c�X׳ї�oV��c:�#V��)]�0�f�����&6؁'��}����U�ȑj���R3m1���~��cF��E҂��W�ȕ�����jM�>__
��0���k��S�<���#D�E���)8����)1wQ�U��4�sPs�K�P��ޗS3��Rr~I