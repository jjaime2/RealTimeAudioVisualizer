-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ssoN3Nr2sF8JoCZSitdN/jn8HGgF3BYrWvs4IuJa/gV7FJXNPK7GtXux+s2B/wdpyLYXs6ZPCBZJ
rLdffnYlCE8rUR7NhJhf3937G+GMV3zG3NuVCWUOpRMcIl+ToOtzUAU5pUcAMRUHDhyALKSr2hR/
zRFVyCtxwoyMrxHI0qltLjewlzq0tn3YaZoPQ2UGi7gro0BHPRYWrJJGGODJZdoR3s+1om60nFko
FMY4cS1Tbx+fY65w54A8kc+4GSCx/R1d8fQFpjBKDCGbBbx8bWpT8ANfSHlnuN9I8boAzO9sIPRv
JYrulHTd1s83lkwsMsyf14TxwyHtieIwSGn8Mw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5296)
`protect data_block
jROuAG/SBsJC49LW0wHHJW4DZAdnxAEzf4yk9TeV00iMDqkULOce8cVy6n//1gTLj1LOY5x4JoSc
l6fpc7wcpVTS3HbRf7s6GOocUv5wM59Bw3P4yCsVgk5H0nHHFOlc99gfyaT5hIPUM+X269XcAHAX
Re5qouKtt8tBSU7n4Dp+ZTRkuUDI/x8EQZJW6R1kzRUEs+QUJDjBSIKIZHcrD1Nzu77YvhJjqV68
d8pg86pd4vkIiKlE/XVhsqqWUKFSFbfyNR6xUGPa/JtE0r6KBHZB4HY4UnEwz2Sd+d7wMwlaLA+C
FBHE9NyFJN8urzlm6acdoDP5Jw0Eua9KPe6dP4B7sZxH0rBhp6Rrsa9V/ChJsCSioFoufTbEDDdw
3TUIbY7JSPhYwZ+uzd9iAYTPzFvMQPSFexoh7PUbrFfao99A1zU1v+uMOvJrhssdxfNAx9uhB8/F
K0wHrstmlhWb/jZWSom5FjKSSWjE2b3IikZ2tVTbn4KAUoMFStBq5UPIebVhVWKcaAhfuHQ28Csv
y5vsQw+ohlJrLQfBlOw31Kqrck5lSoMv4eKSaWAi/rTyYuGIPVJxY+G7IzVjZix+iZyPYUS5i+Ez
o1cvIX0ddbEdOFb4HyHTktAY6FSBtrSWWc1iG61Lh8TcPttal4uIN6GzvN6vv8EfAqWbUAELUlr7
+ZQO93E0anmdLDqdcI8Jzp8OlOk9Jp6s6QGrlOmT6UgCFRFHoSOlCnpgsQxUaOw58dEs2N1WUeEn
lr5cgYHkDitJH7YJWXK3ktu59c5VIaoH2UE6ncEMhtiG6pHS0rkrYiPHfo9VxBoTLuCpgg13qSXR
4d+wsbIq+AfWg5qjLCYON5rYwVLa7fgskhGkEomiuIszUwXZyPdsAfiAlGFaRDqNddNUlSJ0DJOq
z+EZKDc3dq3mdD+7rseRdbE6itvMa0+OeblKdsh/LhWba5z1/MAY0g3LOOYm3xxUoKCkFfF5Rrr/
tarV4vIm5WvCTNFGCcvtIvF3/QB2pRaCcBv2O8IoZuNatM30e6e5DdGKKgfNngITu5KyzgKQwoab
tp1pixn1lKTKQ/Mu45eMH2JkfNOMrph+6dnL3vy8kJiVB6AJLJiRinCAiE9MY1tJJaUOFLmX+Bgl
rWmnIR6E96me1Qm9k/idjtmMzUXCCY2KccSgt1O+5JxfBmO+dLtLRGL9zd3qqv7jWU+aNoRF+DyM
R7o/YcBmfOVCIEY6o4jJ4BV4PbHJA4CBPfRIsJWTvobthhl7d8v4Rkq+MJT0E15JCM0jzrGUdGfB
y2BOUaV5DCMWZHzzr6Od9GdO/Xc5eUsdZ00JQKI/dS2PAXOsNj0TPTGtJTeIMNjy7L/9fvU8I6gz
EwbQWe/0+yQiZSf0k1HL8s3MYCk/OL6/4X6ro3/BvFMfqsqjSEtaeTs/E1FPMLw9M+ZB3pYj0aTt
a2jfgEg/gDWObkkifBjcZnooE2xLlhP4v6jxRrQyIeSmKEgt/uz6HD/reXOT+P8fvHZIUk9fVUlw
oCPthvcBt6JlCmq8yg329CtILLjyPDYrHnv64urff6gVr5OSNGFIq9okYZli2liVqobshnNEsAcm
YPst1mMK3f2o/AgBVH6joLx+26oe/soULgSEwurzh9c05zARtm9JYI/jeG25ngGaAMQZHZTwJ6oH
AYuwet4E5cemQHRJH/Ty0xkI556ICr12No7UYLmyYWgfr7oQ74P4SShk7HkrmKocEI48tLaDBEtW
soBzzxf4OzGrV1dVIuQmvqwdsJpaWressw5CTYDaUiDekuhdxxiAYz24e6bEX4powNJhbGH/nlVv
9XZkxNudYr7GwH4MUX2Y2HGgAat9bEIK3l68LIQDplYfJtJK0iCtN/DsUYmD2BeVx8mZuu1g4++X
wosNCuxZB235LGBTM1sdbblVfmVtYP+8NGd5z2MykXMfgiPawzNGQI111gj6Xyhh1VUnnV0j8n/1
+z3fkffEzPlwPynM/01LKlL74MQATETQHiXbivFYwgTkUZd+ZJQD2nHjZeSZKXj4aGqjPv/tkUBx
JdbzT4jqcvlHuiJJWMinK19NJxR8vrACkOnuqg4/61zSiZHCqvjZaykRITyP6MneVMPlVmuBjX0U
cxkfSP9z0yroVtzxSBcoC6CMlumHdK+9xf+pW23ACFtJ1hBqOAmmArsV0pCDf6KGmXDC0qYsnfqJ
Y0Q962IL26d1VKpRRbZhrBVZZHmmU10tlYZwi3blsiUs8T5jBLC0MXvHzCsGq0vqpvP/45sMt07t
9PKW1lBzfC//OglbwbGHwBfF4vLJ4lTTbtqrkQyJwL3BKHjYEYUphm7GNvmzcfIUlEsBqOZDh6qF
V4PNWxIhZYZ2eKATGmxE4QvmQVjN8VO5ijGv7YelR0taxRQYxXN85qIvRMgRYm2pjIyhkp5/EAnK
fOiZfM/qsa70FB1gqXwdK2cTtPm1NMxy07ITswWcxv5SBE/4jWyiDwxjhI0RQB2CoaN+GRO7xcX2
3mX/t4WIgKwtEQk/nhmSgm7cfLldJTJx/BIJAnku7Jyd7Nhwx0avq7b6nthaE0gPQTbvT6V2MeKT
3atgAivvS3svBvuuJkOzQwsvb0CvVDlcYyvxuVPpohl3fbFGcM6Z6cNIuoiB1Nh0pQA2IScYkhvp
iYDj2D5l+o8O82hyfMs5+Fl7YtslN0WiOJw2MC0ordk3WlTOS/QGqEH8O1eS3XtYxPpC+/GXZIQa
U0ieocn9ICYC7eE6INJa7WNKcEiTJwyUfFFX3dt8FIPpIHSYrbc+L4QrjA1VGR6nyxTULEFXsnAU
fb7vzrH6RuXCnH5EWZxfLzGSmATgq47TSic59kFM7Ybn6o405nzYDkQpK2oYJVzVv6Lc+2pm39Dk
gqiiuuVFTe5O0Re4ZQUBS7/YIcn8TNMl4zT/Fl2vA2GlYrpXiw2DfSnqwkpPlaNpdvZQwVM/WJaX
zRMRNB9tMp3dH7vzpbvKR7Or+54hXfAe23uS+9n1XpLsOJV1zlKjVI8QJ902hGMzsFZR+6Q8MzXc
q9T7KSGxUv8AvTdRvzZzSXl/BzHoKYuGjiQq4nywuowl+rC76mYeA3avqIJQgd/zE9s4NQqI+0zz
+DQPnEAo3kqFfaWILwKc+DmxDY6K4TvenEFf/xwPHp5RaOAEdu2PCfMJJAAucBlqbu8cjRYBEX3h
HP4cfJF15Xy5ryNPs34XXn9PwhjEsZ8o3yh9V53WnIquvTTwUVlpbfaXPDmYwM0qsR1wD3AtMokP
kpOKl/xoaBic370OZaFWGX908vxgtxxp6MS9/3TnepSyUNtU6fsD0MmAfCyR0ATqmggoEt+MXg9e
0g/BTUgaiwo31amOZf5tEv2Ytngv+32MuyDIPf7f1WWN/M46E6BZfF3xhltTu5bf8CAkqZdPFzv+
85lqHqAHsEkMSFcQpK/QdvXtvy4AS/BOUtg3wSsacig+YjyK4ZgnBxU9Pw7fRsy5DApY/sfEtKfI
zM+zsDt9ANbihWtSf/W5ohZE7ABV9eYfPDbh26e0aihI3n4Ej2b71yUyKJ3cSL27e+ozHdjPHGSd
htlYMWbUmmZsWkTiAYJO9hBCF73QT3VDFxtOiDRIh5RxnzQcHEt+s9JiOiomZEUmkI89N4R9180Q
R/Rj48K6XTq2T6Ou54q/ukpawjjoftbmOOgHg6YppjnTEGdTMAOCYISEPu9MFFg28LncjSUCJUnN
rHJfnY+2amh/0xhhLULaEhDHpWZXMTC0h9k8KuThiRkWZ6VwAstf887/xbvT8zm7hZGr7/JHOLTW
zJejzGH4LHaYRDP+rv/yK2JyqRGMCvqJhctd1ver/PxP4zPsGZKpU5z8Cbe4kTGUlcGOIgCErqwD
ihpdaNzzBZLf1dstsD1ehjZl+9qqXwZtDDuCAyaTaHf+4rvcexCTQUMNell1fWgUQggvpZ2GPQcz
4XKOrrz2Hu5lgP+TBYwIoxndPSfgQcweOOkNi4NS9wL7y4NoyUcSQq/6ApgMsxz1irlQsdxRJph0
viaoUif7sn0kuTbufGK0DQmjc9jUAkh/vbe/Z7NtTUqK2i4xWUVWASnpI3UstzVBniggYwvpChAm
CBG3BOAvGRZ2/7SXYRHr9lxJT6/Sv6cvWAisVmTk77z1RsMQKHUor/efcJFlE0L17QECOD1iOtQB
bWIcWLorJtjtcTL2eXPmUx2tUXm7oR1BhR22+rTBhnjiIQal3oDjfqSkmaUroA6OsOahmpzGGjQ8
/ItFwcZh5mduBbYQ6uSs86/S4Klpnu+sOdSWBvFyx1JBeocDcoktwAajTdmAwrNfY0IpY3/alicP
GNUtrRe6qZt2NrmRrL9iUjNTtdqJZe3edu4p2QQIQSRlbWctb8XFtulq7iyALmXpYSDUdEfJ7h1M
TjV8UQH/jrOAZT+uV3A/jsV2wcCGT8cEgSHDXvklGZa24To2eSj27Qo6HDWNj3dLhzCsl6aHDo2y
C7Gi3s7yQ/GwJYZLv4pks6xW4v1S7au5//ixQcjrp+9HmzrurvJcDxzl5xqra7f8NGJaxQN99z/3
H6B4lhRtzRSCFgV4T2yVdQeFP3JLfKrcL8OpW44pBIFLbxP3vWKS65sCsW3jxzXYz11SJ2mFJeTJ
yDPwoMXNU922k8rTrtwMHg+Mk1/aOPB46op3sh0ctaWNGV1YoaO2ft57hWEhDPQO+4iH1N0xDOmr
yoQwwN+M5Sceh9FPv9QbGfqBkES4yKDr2dpSE8LwHLxGm68V+jSRTYaG4PDEADp0vxeh37YKaHB5
ZLEcQKkgIpvQpz2iVnyAyxdQstsLXM++/FgtcN75PNkgs0W7EMqlwmAqbdfwdeM1o1ALJqZv9UTC
gTnoiEA4xmkYAInE29V6e1Uf72G1DivZLauxSHXPbd0kMBSyOK21xmDSQBMkq2iPG5hKxLu9chr+
h/N3XcjJv76vP/POcTHhVBcqTS3tj0UM1ZLmDscII8i8p5XycpiiRC/Qwg2jU94wu/SBWQ6AVs0O
N2lRdhuCOJShRtvSt0bYKPUCBrvFX6Hj9H4AtonEEovCV7UywcteYPm4eQGJw6zMZJUv5MY0tscf
a/d66R+2b5wYA5JHQ/C8kOYI8TtTR44sJGGd+7uLcB2ccAp80fbCCbdg30XOmS/tngE9z9bMSglz
7rUa7vxfnFqxyb9jon/+AGVZXuA9ut9mUbTR2snCc0BFBuMWTnQgfoGfEt5bEkdfIHA4zsZPtQlS
Y8Fam9WPQVt/4jruEzynuL8FOadHA+NG0pp2+6ERVaV05W1Ux8IapUvv3Hv/Xo6NHFjNhjmsHTua
IC9pQxf3iYQsXvR2rL/+kRUj+vW2NCYw5cbP16WmVsn1HE6zZnQOr5KdcULPiNbnEhAPzHtmPQo4
Z/xyELbTnb20L9Vg9XOpYODsJhb+DxlzHpQOt3mUqxABSt+tFujDDP/x0/lHshyGhkTGJepqp1xD
i5Mri9D5kjPJ9N78M5XG/VthIxeRx7wj/dCWohwVpXtAwz3wbxl2EjUkiVJONFOHHNGTh1V1s/U8
l1peuGfwnWT0mvEvnW+UmpJLQoU8VnnAjB0ghutdCYivDAoo0bcgoJkKlAb/hkX8//0k1z5JfaPO
EPQAGIVAhSiBCbMZoWez24jIvvR3CpYRgTuGdg5Vmul5oX2kWb/XB6itPxEWSezisEs9h4lM9Kup
49xYbAjWgXGBLR0AtW7rzoB/Yh0lejQwrxin+zLxoV1F4NKhU5jGlqB/bMoXU7fa//rx+lcXBmd8
rx2JPZms7KLarCQ3tHeNcJl3Q3dd/ydS6XSDMzj8Phfj3AqBdGThmgscwxQKnHMCmKfNb/k47doU
dEfG+CM9qNj1+b/O0n1oVZT+9vcRWcJQuAXhlrD0aC1oNVB9as0PdLIkFrPu1vu8MeuZdZKmHf2k
4bu0d1bWOdAX4r/uCgdcRxVBvRSSkvTStVKxzDR7ZJnjzjR5uZr3BE4g/ysyKYxF2u3qgS/JSV++
Dbe0NZOrslcQ4OEJeGk6m7wE1WOEGB5SYHDpMUH9hpWi3vyYMFuqBEAeP6koSAF6j8AhJ2VGXQWE
lE9bspu0v4J2x+Lyl/qBRUJDAI28lw85/6JVIJeMW8k4Yqsn6guAsoNAro8iLA3vqTH0ReXaiSta
c7ZdDDEftn9Ze0yy+Lx6fxOTdjJetG36YroltlOkPU7BlbZ8ZsxyE9c3+EDx/xlIlx9rBt39v2HS
OqO42rmfkrU8gF9rFcr/x4dqiQGA1SmZyqolc9/f89qlJpULpPUPWGftBgJs9aUiyGH27fNiAi1e
j4AO7/gW6Pw7bR4y3fMAykkL/mNH62zA+Z0W+14V/WCJMuddwg3DA3G/vmtmfWP39/ONm2k/oNbl
fIW/5+5uO0RxTJ++PsuN6SAEzftSqaeLc1gOPywAJKItjQg6FwYfoct0clbYHTmOCw1CDESt8BRf
JJBWBXbkqZ5EvAdDSYdLqbb4yCz5QcvHhOdORttB+hsl2k/U2jprlGcdp5/4es+7sCL1LybwKnD1
01dvhrz2RhY+SeZDfR90zLtNlzY87hqK2lEt2FCY75vss/pYlx/ouR9GvOcB5Y8wH9tJ+UkT3EtA
5+W8LAz7BXIh2zeCXI4mGeGcD1DGcV2Mb16O3L29p/2euliaFlaJMJFbsuCKrX2u6Tnb09rdBlBC
Gl6mR2mS+2Xhd+Ygqn3AmkjkLkqF/n+abLJDyuG/9m8/oz3ShENfQHyVuGg+Qcvd8YdpbhFkjgya
xerFfgzePJZCeCMazmqY3ioiuNkHNArtpEXmTsItdsllgxTlQI+J0rRRrx55FacHfQy/gfdbKFsO
umUMfhH3p5BggJfLV9rVn+1o5oNQ8kJ/0ouzvygaSkORhmB182gtEcjV3X6hQCsRnvfjLutxzK1F
HtA1bZXJtUIi7eDGgGg2vcG0fwyh60d8yVQdJq5cFgbBaVo5uGH2iifoNrbIa0DUulKx+WDTN2u7
mKNJqbTUGphbR3PnOIClAP66xG3QCezpiBXSqHDyKjqVVGPUPaB1MHo2djMaFzHoSeYjwQ==
`protect end_protected
