��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#��R�C(>�-|+����J;���5ǔ8#.5Ⱥ�`0���Ny,�iOK�պih�W���?$���!��p�n�d�v�O ��E��C��V͐+@�v#z��O-ћ)��[����Bۙf����wy=�3Q�?.��+!�E�jJ$)^P��7J6~�>#�xx}~ )!�p���-ؓ����劊@ �0\�\�V���4�-�X}c��L�YEw�`�4%:���4i�+��Oň{�����O��zFI0�xS%�m�)�o�M�R!j�nS��&���h�p16��C��˹��� �T3�] �5��0����j����E7��T�����=����4$�X�oB�M��x�;ܢ>�33r������,/�{���^�t$x�69��{���t��_�3�B��U~c$�����B��V��g�ȿđY8�餼~���q�Ř���E�j���>)�����@���{���[r ��0�ޞw��W��z�A.��^}��TC#�6O洂0���9	N��Lu�&�C�N��|�y�zդ�1�(&I=����
�����]]�]m����wk~�o��XT /�w"����%�Z�����o��oA-ށ�q/{�	����%:��l��/#X��O,���IM��6�c �+��}Kl*�
����D�\�;�)������`�r*4/�F#9���mS".fN5��䪷������WVo��@2�Qn%� ���K�ϒ9�ŠP���J���ўT���訩v�=jIV���lC:�����[|�?������	�=D�$4^e^1�����=�TI&L� <��|]{�N��5��b&��>�~�0�f��E"=����KA,M�|;Sl�դB��|'vU.�{6tvxp|&7T8��)y�q�D瞙s�{/���[�@y99��fg���$��A��R&"t���Ë�T5y:����JL3�P�Vd�e������/c~�a"},Y:��-���od��ѕ�])�B��K�U�?��P�/����^w YN�8#�ϸ۽�q�XSu1fG��1���9!�U���կ*:/�h�jO��� �5�/��c���aS�G	�n�����(�L���{�K��W_�~S�m����M���3�����f2*��l�7e����}�^{����v�3����7�&�3��ۈ����CM$��!A��4h#��zq`����kF��[Q��@R��/�u���NAb$��Ŕ���!͚^�Ҥ��Ȼ\Qk��cźЯ����!���Į}&�i��`�Lr��=�dLa�52�[F��ݬ�ɑ��웊̖�}ERo!�T(��G�?�#�tU����Ʋo���c�k�:͸�kWɱ4S���s��%��������,X��+s�����5j������`��K�#�D�3�|�jA��i2^͌��ę��7�h����ydf����>3��Ż����]d&4��^)'�6!��R��)�����@Xy���D�4G<�p�̿�A*��v�Up ���೴�g8������5�rʯ_��k�Q�G�k
�/�DZI��
w^3F��l�:=x�4�`�ucG�ؗޓ�Q�5FB��7#�}J�q���!�0���#)h4����K�^?\.���ZB�� ���DiS����������,pqD!�Gv��c�f��y��.Ĵ������<m7���1�p$X��g���ѤP�����܊��vQ��i}"�,�%ö��g�G1_C@CNU�`�&!��������W<3�r$�=2X˼�ł�'qzI��
�� 
X��'הT~�-G�y�y�C}E�ӀzB���3'��_�(
Ʒnŵ�=�8��R�-+�'+����%6��� B���1��c:S��EW�U����Z" �J���$��A�S��P9ʕ's��ܜ���h#..�QC� �Gx��� \8�[�f<K����?�ev~b|���R�wy]��њ���d������<��Į��9�zT*M�߾~����0j�������ud �]g��ۊ��qq���N �G(���n!��F�Rz!��g]
a����T�uu�!_��8M�k-�J#̘�=���-�Ӌ�صq�G�/5K�=�7�md����b 8\���AӠ8�ϓv?�ߜ}n/C19x��pJA>oQ2���Ttd+ĸ�"����^��-�[�Asl<&�"Ted!�s�IL%T/*b�ϯ�1s�� 
��!]��1�_�j������5|e?u��Z�Bƅ�.�CV��_S̡8%�{��au�|<A�1��ӶM�7�0� � �ޔ�`rAܸee ͪ6A��l1^eqKU�ὒ"7���w}���Bl����U�C��+��M�P]��|f��l?����}�-��u�fu����e�A��C���.�-g*9�ᐽ��K	�;���f�S��ȶ9��U�tN��c�(6%V#���/7S��R���D*�!n�{M�У�ך|�S_m�Ǵ���6�ޤ\�W����/�tJ��������|�,��rX�{mh3�R)�eK�f!���f�%R�X|5��T��7�6��|�vqK2�xW�	�㹫?�4��f���g	�����آ�\~bv}:B���A�=�9����E�O#l�&���V��u=Y[S�d��<�R��y�<���<�W���n�g#g�XNg�^l�C	���6 �:���zW�;���`�(��&a4oƧ����7簨����<""4i's���"l�%����ԃ�T������̼@�j����h B�6�i�*tv�K�5CU��Uj�U�޳ ]���&1�,3�q�ϕq%eç��!�8P�w�<|W˱$�V#�
R6�}��Z��c	��Ef#6/k:�#�oNq?pZ>���� wҙ
G�6�9@+���p����zS��a٘�:�2b3 �P��,/�i,��e ,H���V ءQ��?�G�=��z]�yK������+�"�Nhh�Pڞ����<T���m��?�/���<���e�]���a�(4�uT��D����o�=����)��mG�q��K��=;���Z;pd�ȹ�xv8��{���y���k��51�S��u��v�g�@c�Lŗ�w4�(?�Kx3 f*{�BHM����6Y�>{�Z�W��)I��(���V0�Zb���s`�՗�Mb�O��A3P 7V@8p�.@����M�O�h=�e6H�z���i��,?Q��x�o�
�����V)�
�������sl������"��������p�jS�1��\
����@@̛)2=N��ƞ�l"�>�7U��U��t�R�V��'h�X���.J*�M�:��R����}�F鈋��U{�2S��&Ș���I��D0�Ǉ��G?*D�v����ǹ���z۷3�b�Gl�&�����`Ʌ����
�u�FI�9k�Q����l�@I¤�.B�w�ꓪ�^�ø���! �)`�Z�����N��ۯs�e �r����C���cNZ�_��o!*`H�Z�<�:������6��Ԙ�B�r��T� ��l�/�hӼCp�%��v�rs�v͝�	�t�T�Qc#R:7�d练���>�w��^WK=�:��L؅
�.�Ů'B%�R7�!��+���g�zo���������q�~��e�\R=tB��B�3#�L]+���H�'�ɗ�q�bA���a#E���g�����M��B%��&z�c&�?���(�Cȷ�/�vd�0k��]-�n5�� P��T�����,�1	��9��$L;�`_�+������NW �3�&*k3~�����h��d<��;��c���2�<u��rxI6������N��R(]}��l;]
�Cb��|�^�^iKI\��1ԔX�0���G�k��L�ls�w2��A�9yWY�9/����*��y�':p� T#�>�E�b&��h�)��M����f�E��)��L��6]��X5F#i���
j�|����_C�G�r?���L{��uӇ�׭�/�t�����mN���3��&��q��d�Xb�6�ai��zw��Og�uo�:�75�Ty����;�1�!���v�IR�q'�>���/!Ϯ�%c�@z}���)-�ݭ/��lnr諷�<��c�٭"�K�f�=����WW���?���r ���`�vJ�[#�<q�Rvώ�_.E`�x��1�]����`C
���S�8*ןf#��ӱ\�^�l��A�9���z����m�m?�����l��8B�]b�"�V�fn�sf{�+�g�,�xS����Q��z��欱���x5��G��#��6z��w)�/�W�`���	`��B@�g�°Rԝ3,>�V �r�7[��K�aan�U���d6�%E
�������Z��"[�y����2��p�bO*�+���V c��~D|؍�M�,�S�Q��l�7X�m��QΫ�� R����\�Øb��_D����N5�I�*~�������C�g����<��bi%�*�e���c�k��&0a-躪\�a,�#]��q�B�}Ium}p[��I��4�";v�T+��|H�m���e�Df�����"�r�uI�?���Q�hc0��~ׯ ����B���ߋ�Q�Tߨ۟Ip��q߃�M�OO�1O�������[�14�'��͗d��K��#]�C%>5m�������`�qu>�Hm ����#�*��<���3ز��:?dիp	q�':N��F�\p$�������:�X$3Kɇ�6p��Đ0�x-�%G���C��
'��ϫ��?����+h����< �V�H2a1�/��[�F$�a�G��W��&a��zx��Dq-�tX(Y㦟e"�~�Gf�Z(����
D��ƚd���^G��F��ꢈL�q�"m��ZE�'=f�/��H�\t�<a7j�]L4A׫퇾~dM�(��1ϔ����f�� Ƒ��9�L<��5-`�m�>`+=���p�:��K>�\��?^L*W��^"�j�?���.��bhU�6�Һo���1(���,����I?c|E�U�|�w���0��^�m�����}TC��D듆;��fG��?�����48�Rz�� ���>��d��~���u�!�5
��^��٧�~����
�;q�'i>�x[ ���Ͼ�t���վf�b�x=2��.�5����j�G
�E\���<��嵱$�/#������҉?Kjª�k�Ah��a�j��T�����b�̕�$Xλ��%��聻��H� �/>e��ŋ�����I��*�kxj�^uH�#O�+�OR �{�9&�y�Bx��xc��d;IZ�]8�����Yc�^^Pi�w_�2E8�!�(4/�E!�*k$mC���7c�&�h|�%?]t�s�������G��ʴ��PY��oN����V���y����
�N�'��^��z�x���vק.��C� ǽ�ȤT�v������^V�(XʾF��y�a��㏱×�X�����"��q��ZԻ'iim���)���W�/��u�Qz�-�H�n��LR�U��E����/�Q��ξ� L��٪q$li�=/��D�|�Y�$b�ϰ���V�}'�90����ע�%�>�3�ڒ1W�.�#Q�m��3-���S:�g��R0�ء�Z�����yϔ����*C焷O