��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	���v�T��_��\�F���&Q�?,�xf���4v�zm^7�o?�π���{�D�t��^�aMH��b��DJ���N���&��	C�Li�|^ce�����itֵ>.&~�J�
m�~v<`��̾��l���K�{5�qZ�[���8�g�`�� ��n:tYK�0<D,؂B`�����o�I�a} ��Q�V|x��~a
��R���M��6��"�2��3��$�U��&�4�\�� I��k0�����;�*�(��y�ҟ���H���7^�l�O�zY\BnƠ^�y~��xT<�ma��ҧ�[�G!�wyz��F��ّ-��`V���y���\6޻�ZNE}a�H[��^Q��6; l�N�8C��`S�3unͧ��T�c��l��ۢ�D����Pq�%ܮ��*����{��莳�EIN@�ȩ��!f��LQ�y߭��a��9�V

�[��o#�QT��G��6�,\JO7��S~0�Z�uٛ@� ��+��87�^1�� 9���8ST�|����6il\��$�H���r�/'�m��;2�=��ɲ��TI�aG#>5/:�3?G����Ϻ����4���X��ü��m�������,И�-5�1Et��5��~��>�ځ�5Z3�7s���CN�毘E�5�05���۽YG�*����=T�V�*��=����TV�.�%_œ�=¥>�OÜ-߉�^�%2g'�sL���c��w= �t*�����x�c�,Eu�m9L�w�^�ˣ�M�Y���T*�n,ʙO� ;�VY�X��W��Pc����f��b���VifQ�n��n!�9�-�y�g~�]�~�;�c�EIP�x5�T.�᜸��
UT|�NEU�x.	�Ro���C�3�����:f�X!�m�~�Z�Pfm�8�صQ݆q�W�㈹�o�lb̭b�����T��W�NI�ei�`����G��pb�%�j%�J2b�؎p��C��o)7�`�`j�-�w5�����8�L̵�ra�b�v[�[.�sJ$fr1E4��;˒ki�$N��s��&ׯ��A}n@q�ܙ*ɧ��nB��E�N��I"d?����9az�= (_�J�uP���B��ePK���Y/���謷P�kJR�֤���9��zU�Q)� ~gH����.�*�Ǫ�V4p(^�F�b�ٖ�AB�#�t��X	���銏�	�٭-%3�a�r�Hr`g��E��j�e�~h#��/+����_�>aR�p�������}Hֽ�����pi�Ɏ����Om�5g�q[ ��y��q���O�\)�SWR��E��:DXH����(�MA�a�}�r����ZiH�6:Z%�i���>±b���i3�O�\��>։���yA@c��&r}�����~
/��U�vT�;��������]K�A]/cM��)����N:ᇴɿx�4� p'젽����ׁ.�J�p�g	o=H̩����Z�7( ���D3l����pM���2gU���|x牝�UUl���V�;!�A�CZL}���ܲĺg��c�wġ���W�s��^��nd��|�&3�G"�z���6����)4�c9n
���g]x�Z��7��-
�X���	���WR���{�3�P��ﭩ�<*�ۄ��q�Qa������ Ol�60Y�XN�%I����f���"�p��8̑չ[�畓���~p1�3̀�a�
!�1`�,7-FL-@-r�z���z�:T~���Q�{1�H���wJ ,�C��ѣ�L�����f1-�[9]%ogFK섾`BM���9��7n��	���E_������!�� ����y_�0 kqZO�O�E�FwQ�^�N��Ā���;� �,�^D��]mS��L`<��dʾ�4�rA"r񯱘��i6 ��8U����M
ѫ���-�@�sy�6Xc4orW��b�}ޅ2D���P
B�S���Ot�v�0�)=M�z��L�x�*�ڲ����ԫ(��^,��\�� w.pUl�\{.9�<f��U�Q^-F�m�a����j]Mp�]���:�|�ixuk�~(O ��R��n��;�'F��M/2]��y?�RL�y����+=}S<5g�s%�.���+^��&T���m��L<��&&��#���TУ㈿*Jn$��#鍺Y|�r'�vb����8ݱSq�5~��4�����\/�ZE/��v�0l�P���[l��b'���N�F����pHK��0�Ӭ���t��0�'J��o����v��QE�$f���爳"���Z
�'� ���f$ru��Rsj��$4�EB�BYW�a-53��C*3�a�N=���z�i����h���/Х�2vPC�I⎧���ߓsQm��C~�w/��;W6;.�aB"ę�ʴ@c���v����,ǈ��I|����<�L��-���*�T��G�\�}����+��NSAa��لF�3��VE�HD*�r"����/.��䍴V ���^q\��� ܶ�;4��5&�}���o�C�o����������` <=�^�ͻ2��D�~�j�ūqB�S�auq�������@r���k�G�{(d��}�I6����yDE�ߚ��%���_@��_��9L{c"���q�v����:��EG�q�z-�MT�I���lM�a��&�tکf�=W��Y>��ȟ�Ue���!�q	$͆Ux<������)��"U6�j����y�r���l��ܠA�>Rb�p���r6����w�J�m��#��܍Xq qVv5�g�OÉ�i�<T�Xӎ2^L�C�5R���>��M��-g�)��%E�дPjfV���r4f0��|l��|�ϮR�����a_>�1� �*%y����ž�@%w��3fꦹ(�>N@���L�/+�����ms?e:B�n(?t3��لR?�T�j�t��7�������k�$�e��s��|�Ko�Q>��.���>��l+�AzB�`<l���������RLoR¯<�g4�WH��)��m���``N���-�j()������G�w	
��ej�M�W����"�^�~+�93��������%�\�9RRS�.�m��:��=��़D�뗾�L]@E�r��7�3m��iU@���t���wL��E�Z�T���
:��80#rk��ͣ���-l�ml���'b W:=�5����~��e�
�
&����3�.�U���W�#���ѡsպ�T]̎D���0�R	xn�K�r8!�<СD�}��F��6N��)k�:syI��ߵ��_R�MM h�D}�7"=�RT��΄O���=��؆H����>���w�&���NC�ٶz�u)M��AVo�uܕ�M�n����؉�8�Qס���@n� 6������uҗ�e�d~��@�� �
NK\��� -�pgI��aZ�Ka��$[ȯ5���-�ܿ[����k�h7�E�i,�	˛���_��"�����P��弃_�T��F��)�sI����~=	Q��*>��nE>wqyy��M�����%���tW&�r`&Q��j��n��H������1Ǝ�8X%���L<�vhEvw��� N	��4m��#S��&R��J砧�{@�q��W%^S�����(S<4R�PL�|vq(-��$��t��S��B$���|�!.�w����]P�fD/\b����t���h��bAR�ۻF�iE3��?�ؼ΂�x��y���̩���ޤ~���1>Fm׳wA] ��"PдN���\L�w����ĵ)�P�����K@<jW�5�||M�"K��s;�4}�KG��6+,q{��n�3�i��1��92�K�� p��S�w�4��-�!�����\a����m E��_@���C��/'Pms��T����_�c�~�[�V"���iT�^o/V�uv��)'v�G���@�C�1%M�k5��x$��7����K�P���@���C���h`I����X��?�L��y;���	c���S���["�Fg�s�O�ސ˞�r|+b	*��.���ϩ�H
\�(3^��C��	��x�@�#�j�e?��S!���̇�/*�d!R�f���Z>���E6�c^/��n9i#�`H3��	c.�Z�Gb7���6�,���Kk���~w���:,Q�@��t�x������!��z���)��D�i*���h&�u`*�z_9՝	V	�/N�k�n�S�_f��^3{7	����w���Gf[)�Q���^�)p����C��e`�='�������|�u=�9B�u��g�̆��H��T�/1n�� cZ8Y��M�j�%���u����5�����y.V��/k_k{�P@O��@�K���J{��a�"�u*�O20\rTK�} ?ɍ��j�����}���p�K+�m��
���Q�\���b��c��;J���7z�wIG�4
�����&����;�k���	�]M�Q���h%ӷ��G�'��+�U+�H�ً�G��O�!����"�)�?b�wdP���Ʊ�=�t��nk>6���	.�:�Y�e�Ko?峗"L�W��L����ޗ��z{<AVٗ��$'n�iZ�[�/mc1@؃��[��S��/^O�����F4����R���\}����Mr��{N1�t��"��>`P�c�ɿ�k��ׯ�EKՇ~aDm���{^o��V��
/V�e�����>��o�9��+��h�7��S`�u?��@���	Dk`�U}|S9����I�Wr�ϡ�Kݮ�w+~G$�����9�	0.g��b�&sNBUM�����=��1<����n�#5��;�i�݆�I�k��y�u�ɣ"R.+����+E�-�����U�o�ϡ0�&�O�ť.��٪78��l�#G�g���Q�0+\�A*�?/�,l+�F���U��s6������Q�}���-��B�/��S�7��\��Tp=>��b�
���K��;��>��)�h�2��`/7\Y/�S�u?ǁnA��o����f�PP��ɯ|�HL�Q�s����