-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fYzqq4ATUt6eQ3zro7ueHWGRc4VQ/e5CntOO34In3LytcgczUefnoo/yOZ2PHkJjqJRU/HltLXGv
tEVKpgFFdsHfPW5wXuSdHoTyqF/Pa+AcG31ZeoYD63/ItJWodTWB66fdPi+3Ten5gqeS+KvrsxKf
vBFflLZZbs+t/ZvuOVwm4S7RAFrmg9XcI7gB9jyrWPNcyZC/4tWBBNu78vjhD/E2tjX/wUR8p1Mh
dgQNgMaGHKoAtz+hDhQ2S8/vwrSxRH4nZb4gRzX5g30LV4xMprCihUtS9EI4Q24RFLkV/ooFarnP
u1luwkWq8hzedLtyCvnEtq3tSFMRkv7e84xfPA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
gsLVZaeJHlCVGMcEmooGO5bLE42BNNmt0zCr1oRZVS9GvQHUqP7wdVsKOgU0HrJJAyJtPmI9p5qp
lkPyVzo1aWPaIZiMCOfZbU8Zp8IkXfSPkm4B5JikrsC6t1NHkdieAM61KHRP6bKY7qSZFzIK1yyT
roVcz5GpuqQ8vu9eUEB8sZDVyw4JE0VuLPkhsEgRdoj9kXjSQpVMVoytU3CDFh5mJRXG7K1CGq/M
DUIhEqyCRpy6O8QtYzmDYraAVsPXWQxcEUV0SxaURDBW6szEo68wkR5O/qcy9zq8vUARCepIA8vx
3XnFTa95cTTeoxxG0RWtpRCmn7eXYh2QxQmkcG4qVfGeK/HtJLHF/1wcVVbxPYkKTcDiOrnrwphT
TVj+K13FhorIzNsSeHVsWcquFPdwuoEwmHZVlJvvxw40/JOsiqm63gOWJo6We0Miv4uxt6GAUM7G
6EYAfcGuhBvhNlaBG+c5gHJwvyO4L26gIQYf4pw60lQXzaiX/COjHZwa3dZww/1053+V9gKS+X9q
mbkm0/jGz/udiZi921r78kdgiYmW4qhhigZwkSZABT0HFbWZkxp2898gbF0QRG8fgjQ/TP8kyvVA
8t1zjdRlexBIVGgmAevNrbYkf9ZAAFIoBhgFffq5XYtGM2hnLCvV29qXpulHABbTPdyeZKfFp155
rM0BZOH/Weae+WUlMR/025pNAwrRVW4XGoAgYjiOypg+MIW4OL97HN6mNQTE2879dBUxBsszNqdx
avjy986p6KA2CEz6dJk+tpVoyVrk7RuXU+Rr06qYZzag+81+dwD0qh8HjgmuK/vk8UkEJYIzKviH
ppHiAo4t92/G9qqG3bJ6wwh+Tma+RpOzB5hc9JoSm5ZovGF8XtuzdMqEtbx23d/QJGlVCGv+H3LO
IHQOEk0mlWzu7NgdR68pIA1nBYpWvHnJ3JSs3jsTkMrcThPFCorBkqFJxLReJlUymL9Zqt8KV1i/
ZmIru20a7/nEElxAHXwk2XKlom+hRDIGZLbs5QXgrrk4FKL5S6oJAnogc9RUFtYiOijKbBapTYVN
TDW6FrmgJJAv0TfqgjWyCzBUGHArxHKQmtBq9Py3TGnQN1a06UFhh/wdYN7lTbZjBvJkNhHi6o77
gAsKf4sU52AMQ+8L9qK+nu0Wk7kL6FnKOrsU4x/IDwSI9cMe2lgytIHuyg0O0BJBUrIvuh+1njiz
Ec/K765UnQXI34yzKYaz1YDmIwJT/fvXHIi/1EfSyVtefYHwb/HQKT3Ke7SOzS4cmdWc+zejRWn0
tDXf/p1k7dPYj+FX3QZTPaDE8B5LpyUN0QsI0dEnTCWRHKrKoi+f1lG71UzbEjWxDiuikIiv4ReV
bRZO/YRly7Jk3JYQ20f75Y7KiKvLg0VU8aQE+Zff6aP6U+/kA/Y86ezlXY/mTWENE7tFkDcrwo5w
EsdzJfsptJmfTxboNv+u6UDXpy103EPkvTvCc7UiwUVWooc7qu1JbgE/xFphCYLgOmBBG3Grbbri
GzD3FPTMhci3MO4mrE+6zTWHrOOexj6sgiqDMYy91vzNlLNhhkh9AsGFYYbeDMshaW1NEfAaRLCg
gMLpw9morK1fhrwQorFyl00JWclUR82yiDcZQVGdTcqUK4OFuD7zx2KIdPs3RakJ8tumSqcQ+/Uj
qFxB7T6CywWLs8L4XYyFTA/zo6FAXTHIPGk32ivZIlhUk5dJE+F/M/Qigb6blM5c75zUnrPrcox0
07j+MFWKrgVDEff6si41G+De9xhrxF2fVWbnZf02xZp06Fa0NrflM5RDnMZ3Hw2g6wE5VNWUVWaC
yv01uYSaXBOuOqEZFc3xE5iHBB79B+MNMxfNslVSuxqqv0lFJ5J+LIlx24PUooY9XOQHD/qWHMJY
3HQNN8Lmuui4MNQn3sbwuVoo5Lmaamv/0aprypksvVAkTlLdUt73l+MvwsEp+jBNRcosiEZTFX3l
sJ0QvwZZBfGZA6QgamS3bHUPb/790WdB4xCuGMOMbm1TkSRc3HK44pqcQcE3lDqMpmB+1O2Q9ELE
YmJAjciKe765IFJQ8pMG/y3ZREU8lqZ3BkJwVvwySI3rdNxEO1MhghNPSr2QISiRSRavvdf/1g9I
0Ee/Wf9ug3ihhkPWFIbc0+7tFLI4rCLYVrEwyBuNtKcuMM2MI7dVeaiuVD1W6v584UXP48BDEE+T
o6+kRwL/H9e7AVVcmjyXV1kFIhjEvdl79tt/zGLZNtLJEYj1HEDBbWsdk21vsAOG3KHCcJvuvi9i
VzVhI+fvq4yOU0zno5llFPXQFkIvj7ImnM8jQkb/nYGs1aCD9908yijN6e3OI1svLsVlfmnIl7XR
HfaEZOqd9vlFeofJH2aW/tBCJUjQOLLVcN6FZHGrk3Kg5GhgbJxafGWXxBQblj4exqmLcp/hnOOl
3hGIdf13dUjzQunrqVund44B3bzE1cGdgw+icKShhCM8U39PJRvZymW6KEeI61vfr6VROEw9omzz
XVsJ9kwut+8mb/ARyFETYFbkTxByB93jG/U03eTKteWFjfYOITlzoUsRDkIg8SHIfvkhQggFFM2o
O2914p1I6TupTuf9e33NXt2RXNQrhobRexiLBD/66ePAdVSx8qGikEEq4jx8D1DqKzqLVqjv1Xrk
8ojvKigaQlCQVVxgVTcGBCjKz2Ko9dMpGOEHF+66nLrEknOviCzDi+eWAP4YTOsHpvSYa/7HfIR/
8TO1u2n2EyhQ11tNEMDK8NEDKueKu7aqSUfcU9+valgSDJJGjwwgWaEJvqH//vmMTSklbGLKy7jq
jXX2pEQR9LBsbhwUOim5rzuw1KgHrcnfRqcIiSzN6Lh9MhOZ0D+cRzAW6hOu2Y2nxOo+6th+nOQJ
xDMK4Ec6aTgnHvQh9Y5cqQBKwIwjQSTRSAq5RJz31sJ+ExS2munirb8HbR41lPltpyFBdA5MTAH+
GfBwOMMGYGCSGhX7J/BUv2+bsOIeiuEmFOO+1FURH4wNbb3C89T7ThH41S/voFqxGPoWLH0pFQ6I
ysnA/T7YwTRK+aaoNSTDoTKOzmEBp+nyf5ix5h/Asj/zZBExJWYXHwojO8K6QPwuHy/l+mCH7xQJ
NuyXdH9V63qS65hCTmHU0FlXRutxsEXe78VY2fy2skMD1io2IMCkM4XI2vcuIdGsli+kloDVliKB
74zRptjHnHbchax/RuVi3yMu3W6fiHq54+xDjim4ZHZ8HQKeoihnsb9Ue4N9WvE9EtylB0BhoFea
6zytRVsUANrbIPCg0V5apjXm2Zslug3SOajGIH6A5GuA+uoJa1lzDcNo5M5aIw/Pc9il9u8ZvpMM
MZxpbrN2z1kBWTJDm0UfACjsNWJGtfdBf0agghNB3E2+9acJsN42O0h6qRfpTdlkc8ITci86YQBh
+h76mcbeOvknVzz6580E9bnezLCHfp6YmFooHH/kld8lThAUGN3kPI2gIAs5M0rnIMoALQgu5XAB
RRtgmBX4AHTYSeCLAJCpYG1fqHdIYZgebq9vI4qBWx0wZuR53YODv7zG+iUlgIBCfvppS+r0I4z1
e8ym5oZOf6ufqv/FJOijiUqxFaI+Hyusfb1T3YQ9PAxMHQovCfSm55rwBW8/BgM0daieiNbIO7m3
TICaR+c5wH+xeJKSCKO0JNlA7J1/oFwOOrqU+kDFoMlQRpjcEI6TrNus63YljbvpwvZ8KZTlua+f
HW4/kWsdqWBDNi+krLr6mUSSzCaVKLn95YxK98T9EIKTPGt9O+3N6QlfkOnitJt5D6CcIjDo+Ra8
1DyrzBr55X1PY7MZBmUap0CaEjICPQJB4TB1mgrocIDpH5DeHLSCJv5c8YkRsk4yiSWPLmu7+Nax
3rYMT+lRTeBAhAey0p+hnNlu3MzElqpcq71pO6Z65PbKy0b1vJtRK9C10RV+zf2AOP/NzFe//q7b
mW2CIXB0PleXKnp9Tc7blTbMpRMfNfcXiKSa3XGFp57b14ZhIfEALgT8NcmSXv5Uf2yGQTAmElbZ
JCv1hMQ5I7jm+6wsrufpSS43ktJYiqdpIM0+qJeC7q3OR56vklMDtzj9EcYgmUoeW572E4MB1RtV
GnZ0XkW8RPMjMEmQCUJvlwVHG5tIe9bnNhzlv/G3x72Ev1hus70ymhpXI/L7HTlJBrItmNBnWnGd
UzmTu0dYcWP83vjqP7gSmR89C4vojj69WBGhD5LOCr0UgZdGGMX/n2xCQnV0mQqLsR90pmgPwOtX
bFiEh7EoInECQmNQWbFMSwoALBIvCDwb5OayWOArbLNLXb3lZ+WLdAxtJOgILWCpMPuIiHPYhduL
NBDvfb5o4H18PFN1V/rqDAG+SRCAC7yVbs29KOlMvZWHxVmAR3AL729HWT029J8Xc6oCHY5HLlzi
taOw1q0uR1Qh3lx5B6IfUz2/wJJz83z7zzyiGTRcCCJJ/lypk3w617s8dyLCAQ8a/nD2ls9VkINO
qt94euOnnVVGiMYh0kcnRCHXbajnp+Jcq+rC5dD/2m5skUd5GLBkzkATF4W7dkBRT+RPkLNuIxiU
FYvEIkS9HD1dT0PSc+XKyExnemgSar8B3uR1vDjY+n/Q/vTzbk6Mq+4nAp1POdSGlIxEN7azqcvQ
gwU6KGZU8O58sVlbANU/UunWzLTv+QPSyz+cMsKEu06InAOvpRwBTXfEydly0eO23w6Zg3Fx4or/
t7UyBm1xktQDbSgIChOoG3LDWuHHGM/hq3LObLYSItPCqbqFYEev9lv4njtZ70Sd0YH+3fiQ6MKT
RH9NM1E9dimGXvZWvi+gVlMBOo/BTkrpux/jZLfngj/wymMWhRgZVXJO0yaZvkdu0me1QvT1Q/58
FR1/eqWYyUsZfJiqnK9HyXynmAlnl46Pi1vmZ++ex9Len86Th0jse8idJyTs3oiTbgxSxFlsRqA6
iDCgfpnsITojRMbI0t35cf0mbibHFu3GsOThEkycbPGYUInE4DzD+x+xYDCizwS2F1fNHEqVYnwz
aDnMJetjL8ExxALYqOlqbxJuak2MAsGFx8ZrzTWK3ldMATFSH9DZDOwRyR+H55ixZpsC8h7aYJZb
UfNe87T7V3L8alzOm3Zlz2aQVY4S4zOVdG+lllYjQxR/GsAgioj4wX633vjpL7niKDDNzSzi6WVa
liiEv/85zI3BpwRLRIVzNyvVVHoNqlv7491wJReTFu/u+QqDdIwgWfmBiOPu0t3G5EzoYuejIbJY
jxvkD3QcUEil5ht6uz3upygRB76wHncyMOudNTqp0wqeV4AVhKjAPxLX1+3Vcjp6FpAFPhmdciZj
BYMPeLFcVnndTch5nbw3fWfnub4zQX80F8BhD7cf0wnU6cRec1yobcjtPHfJW0qGoYqGG8stoRi/
7qrHOGQRQJhqkXDHVYv8cgeVnkZb3OdllHjK3Zu2IN24jySGHRm6sXH6r26biT4eE043vRVOyT8m
WnW4mO69yVv/8kWgRAD5V7nGUXSfuupRy8CHH4NgNT03e73xiWeoRanvDHxq/lBSXIO7mImsCcSX
hwqALhMRZfbIbwSpj5/vV2V+8YXNcYyG8K5VDzWo1WwS/MsPggtq03kMcoVNhfTlthrIvFD5/zap
XfWUrKa/r/f60MUw7l0dFchYYNSs96D45pmUywYoiaIAuGrMUtQMDXMpPTeycpH9urKVoHNtz042
PWPcMtDemnb4xDPmNuXrzo0XjUXDdKQLUKhgaNlXra1YPGR6q66mGQBGKtqpWqp51MBO25NwBduT
teQoiDZKLUhqxVT/ckckW8S54sXlglsszaADEWEWKqbVgWRFZqPf+I9Ralu0ZwE/cEnx8tUmuTW4
uwLFuU+rXEPYLEXdVwnrctyF1ycVhiRGRDxyJhgw7QyT016rlMFWHOJUGY/MTcgXbyYQlIgOQgCn
SytDGFmDLhjv/62kaZp37z9690epZ68x2lRVPMhhl2OeMCy1JSmCh9XAEo3QAZblQmrR483L25+E
eDviXJyaIJzZ/MN4OkL8UEsgABSw6oqMs30Vr4gZX1HspCuhYZjKI6iuvSwbqB3Y3fcUR0j3srMR
TwBjJF1HeUdy1VU05RNqJLwOmTtEyQX7UyPK1xmaqJ2IDNZ1wM+guqvxvlRitfqCzR7TPOABh2U5
wK189krFaHbk89HiWp2Wvl2T/iYLdqT0IlvJ3mz4d5gjT1ZI01sBM0mI3qtxDJ7S7FvnWfieVGJ4
S3uGtHSlQDUj1l00vWpmKFHRpPuQJUzAXDYbn4sU+KEy5zEunI4Og946v9HDmLvulahAOljIX0n3
cS3K8y3MquOSOUz430M/fOoXTwyW+IkYENVLt7exILfEAqVkz0Ds79pIEX+TxHbj35iGBBoNQS5H
A+0nG7y0VVM8Mm+CQV3Ltgm/iodrxohLU7XmONkyr5hOzERpF0zR3QBbn8mRdSj/kXla7tRYzvz5
mvIwYiQNoRhCASxErE4U/6lEPF6loW1cSBRkK9wKRxz04wgOGeOSuOyRXX98s+H2Q+j2eN6A2jHv
QPJ49eKR48afGXGmAUW1MAw8u6mgpUJ4udQicynj0z+ZPtLaQmplCpamMwpqzlJeRS9N9HaoWAz4
IAQGBPvD7H4m24g3kh6Q8CGE2aevymGTpNrmCGsVcWXqIfjV8ldVyYobXIstUGMcvoZx34ffn+sZ
9Aktdbg0ZNN836+RMupB4Y1WIgshCKCHEsA4SYAscy65dVXypW6xlgOTvrvyTY0gsJlsL/j8U64Z
ZVUmUu4owj/HCuARAqaQztwyE5lI95lWoSt9XC45sngLNxTaSQ19i3tIro9OaJPEPpOH5XH3UrSR
5F5Vj8jLhOD0m0SH61QVIwqvx+ALCEKcCSEFcOF59f1ZtzcyHPBPE+h5nefjMKqmp6PenLhoSmNc
EIkUYjERCP3ilGb/UBG15fcQaJu/xdIzunzVbG+qdh/nH7FT+oE2ATC8UDtI2jItLIIZQ1HwKBFH
uf3BTDrvgspgwPjsd2rdA36G++rkmt3uUODlxVd255MM3cbF84vvd0kQmhKwdlzLB3JhThpeNQEs
Xkljepn4sRFRdwf9Oi3RZzXbdBxQHXkTmYmLbq+pEsS+BsgLP4DlTx2BjuU+yIq4T6rnpJ6QyjKv
vQ8VMrdrFMkaxliJ4dyNyIj/YL6kqZ43zPVnoeB6JjUSHHEETqsBlgtmViI/8UJAEYVQ4zgEbAPQ
wA/KOQp/1j2p6emLNkpomjpZPVpn1TCf+M5B1m23tYb/0X/3hX2mkN8z4mVTmdqBw6xJDz4wGBcJ
j6K+Gcg7dvwdGhHf8BkbebwcEsXnPM9k/1oSfGV6fyrczbFw8Miafd0lFPtohFSO6d3/1qlUDgAV
FEHu6VcwU2GZ8z5HRGPPB0HtB63yMAc1VDIJrUk/Lzq/7E5cZlyoQaK8c4uQSHbOjfIZYUSWHdSJ
VzJdhLvEfe6zxEKDz6iHblVkBZdGJZ4S9E3SDRwDrAf2epvG37i+alEBVNpQQRYS/SQ06AbllDMG
c9dSk+dFB1A2+AAaKvXCsj2jzs3sk1gi85oO4AEmbDWqkXvnSGwj1UPcpHI0CV9v9iA0LAwv/K7p
iw8zwqmmcGAUs/bTXkyS5R6p5qOylNHGl2U0R/7X2VOHB+4kC5CkIIelHMrfXW2ZIJ7mGIq7XzFD
Vln+wb9C2Nd3k9VAvS2OaOc8Hr62qUipUKdIB/njhrC2VMC6zDKJzWfur2gnSRaOTvG66IYt7MpG
ZLjuSG9fStKCviTo/f8TgrbMckl0hNratBn94yy6qHkrsiP+Zk7W2P89gYFi0mRbGZQa0Ql6nLhk
FCG0I+62J2qPUlruLLV4JlEUas1b8U6KeODP22McBDYFkh2vnj6EaNtUC+EXgoGZJJ0DfH0XsvX/
SsF65Z3ipM4Il/T/BRD+mePLbCBgsqRo/aMXzyFfKDu6coNIFLE+gxuLKn7PIS2ZTN6qehDw8suC
MeUmXlldi1uqva8csExat4m5MDbvRe/ur8EICG+y/O99TsTOPlUxOTYqMYK7V7IL/tt7dA9DBTKc
HVYa1dKzyL3CgToXNF0hTCy+qbzsl518jkoeI0avtP9m1UjishsFlXrXHiNY87EAwVG1GoxIlqYB
ocme4pT2bUXhSJ85z2IUpIxtloPHahh34pLk1wFOKYe/kFb7aikzN8XTEXVVhhLk+1pENDkSTaAP
ETDBQdAi+vMJy011UfIjIcWmiJM1H3fKUW8i7E3DkQyMOkmKx53GdTOe8/JlA/WOBxKoAs6tA1W4
YYjrxJ6ylAr4w7dAX/rDin0mnH8yN/n3Yey77w7T3zdn3zwjdRteKF+96e0V+15ib4CtG6H6pQnr
/6t8xWzZ9m6ph2TC6lwGGPqJ67PTCa2NTzzN8D/RF0AXpViUhg6c9mai0VpyR8smhUeJN8mhinv2
1tb7XUo9FqjOJGyd+gkQvuzXAzNko/EPMVYnZdO5qxEiMHhCx6uzRd2XDvjXGsKhT3hIs8Pnfulw
rLJQ8WudKI3cc7IsW8Qh2sOec7qid/fKPpkSrMyJiIrAupxYPJQ7/QYdiI7dYHFJjLC8Go+VN/Lg
5k02pwbWg1xEAKyFXy92HGMb8anexsRFi5ziTkqs9Cz1vbf8EryaSn+hnHlI1yH3pUvg/frR9m9s
I5pHWAtNfnOveBgwzIx431uOY5zuzKXyFslLsVPw2VYDSORFM6QunNucR2hYFADHA+vl3V5gLs+h
KcZsldT0D4KFnJkTvhJmg2dkFcrymMf45a1F966u8xKkJXfIMqObzfIG1MaaOycXsM/I73ovRCHz
1yj3Ooqvs4dlvipZ/fhNmTnKFSp0oTghLBP9+fpmChQQ63qjF+skOlQGYuaf5Gmv8jgenSPkgPPa
wx+Xocsp+nSbXh4EBo1D0+FweDn7+Z5jDs3EmSGkMkTlMSBBfiEAGY3zd01JAz/+vepieH+tUSPJ
pDdu3ZXR4iyjYurAlf29Ll3yGs5n1gkMgkG8QoXlPHNiCq/gH1XBm0DMwni3e8UASMe0Mr6ewxOD
itQwukBmM6+P4369px9Z0BZkcLPIEGGDNvFuXYijElzZPQjrsXAImKrumX1d8RECtqse5C+dm6c2
JkltFl8/dJQcL53mUm+/MBYRIcTFzZuaKuKnIe7U+9RQho1hvSsPK1XfkDPMuPa4uauvg8m2//Kr
6TmsN6AOPM3mTLpX+Qq7GPMBRhb4juxxGmhN+FPeyT6VCWudmdr8MAjmhb7MuRAwg35pBhhEz1JP
MD9jQ+NgbbXg/dgotVsgNJ0A8I9ComX05pp7LHSkkn0+3wugQbJQeSjf8UY3qnbd8WlXjXL0qzC7
rLrasmI/CUx1p6zjhqRzQumekDMedWvaRe0Mgs5RzamLh342yYdudAOTHvqYuiCtzDFnif4XlO+M
S6jb8ZAIEu5Xay2hHmh4HYE/pJQjtaDoqLtgDgPA80OJzCproSQPHxRQUDG+9mo9X6zBQVI0sHdP
b/R7NTf/Pm/4jU311/3GAcyzeC0gittJEGNgIEpwCPtZo8qwNU78vUKipygaHB34denmr2IgX09+
OP0o4c47L4/QeSaoe6W8zVZS26vQiabp7x1JnthMlYu7W/177caIlO36iXOvum2ylthRD/LQW3sz
2hFX0Dm6NqWADr6CCLLEb02YaqeuMiECxLNX0BZ/TvKH+D2PUr6Qd+kQZimNgdyAnB4XAkyOUquW
6D/eBPI+jTrr7iu98r8GAjvIQh9a20NP+zn/MSFQ1rG/+SYJt4DJ2rRNMsZRsqTvg+W4u6BUGMcN
y8JpPSfqK+OmDDhfUchHJ1NiDi3rxsEk0Z/skty+YrseyqHaE22gRctTV4w7vGQ/0Pt6ifZ4S09n
Qzr9J5xqQCfuhYOTJqcS9fb0qYikFbQWGIsICKV0fUB+yM4EsiThw4nX5zUihSCUgebS9V0LKOO7
uxMJLEsbY3YzkdNJfkn6YX7CeiouQvUl+svDhTESyYg+LHYCMIB8zeXbkIfIAXxTCKbUPJEHT+iu
yrEgEcMJLKkRbVCiF9mWovM6NtF3mjfoyClf37Z78Ru7sY/FEJpfa+x4nzGBUhqOH6JC0mU6naQf
YJgnycgMxBOCc3sgpPVn3n68tMH20oTh9DFw6ptS3aCCJTsP7Layw/06ruj+OAp8PQgDCkurOjA5
HC22iopbQzXOfMfMU3W+ecaZ4N2JY3AdCKXDu7G5zTYAgjeI9iOk3CrNllMJzsUbF5COt51aKgWd
WCWatoK7Gu/X5fxBi9DKm5/3ysX+9p1SPJaZwOLSJ5jdHbMnkgyH9zk7GLOzJPIcJaMqZHgs64tp
I2d4BVZpHclIr4RfF2RVkQ0UHKDacHFnj+OwTcWPOrpZ9E0pFhV9VWLb4Yvbh19/zV9FuD5Rs43j
OXSrUwBImmfONlQXBAGpEzkVgxSIrTkPjkekVroEVjPB7VmQ29YFMKzK4QmCoU60dIbeJ/8cJ1qm
VBoEp3CQGqUgnvj0PRr5w81TOFaOkcXcLfD9YrgplfMWxGbNRNq8ZsyXutJuqXJmWkV5haTAqmjx
olOtuZD0VkfPqjK6zxjEh6CytvaDhW3bs6uZzSuIu/6yz5+KYmC+AP3FVDwetmx+2ryUL0BvODZr
LCvNZDgvdKS6LYTEn+zZPP7DLF+IWUEVYgwD/r782k3EcrxDmBcwaqT5Z5ioefkeiHxSzb6nxUQE
e0I+0aIiJRhL71SZ6Mxg9IBPEMexPiS5gHw/baGCjN8i4S+dZZFwCiPuFOdymbElY8jUnIv4Keyd
MF0U5rbhc5vXDxjhRFogIgZWO8NoLOvLerjwCTpIv0L8vxW85lugascdkbcg8n7ERQ5JhC1avu20
oLDnEda7Wp8la2NpK8Endg+bjV5TDEVy3htLM/AlOfDA+Ikvmh6/cnQ+V50CZ7zvNI1jBKa0kq1U
HYeXWzgH5dZA2RVCGEUNO0voMqfEFu+eMUWYqql0ChD8b7RKFHjqJ8zzBYp/saB3bBu7mMMuHZLq
WrInClpA6pe4vwDm3Z4KlEu/mhcSYzJZmNuNhjjIy1ZruniyTwdS0qU9i3VQf1Yru3SnHa879I0g
WK56tLR39+qiOah09YQbA1Jzd/Ib74lqRgmCFOXx1N0ksMw/KYzn6XlIMDrz8zmZhFNT2Z3syWI9
gOLz8LqWP8EgBaHQ0rFVeBHbXSPeWpVqaFBnbyJCBk5Bx7g6RxLxpgqquvdqLGCcPHEW8ZTZiVel
xewhokKoUAYJH6YYu5KA6Q6whLDsdzM0To6RrsACsgbKlfI0Thsjcl5D2W2x7gcv4pQLAzYriqnP
ImwhTt50e9vek+Qk4QUeTDoO2LC6pRjYnD8uT9dI0kPHUVW2mVaL/tQZC00pwbH4/pqs+bWJFM2s
qp13lQAWJ+a270i8bX5Ce7Pgx6Lafzu8y11R7Obvd7frNeUR7Yn5vVC2p7OwcThAtfXyapQ2EQrl
28N66RJ+ZUPpN3mKahXYrvaWIntsEomBi5vVXXLTLXRfCsY42ugk3M9zeZlsQT/jGo128Lg+IvNX
Ff/bymcDsQb+9GCJ33unkZ1a+swB/N6iBXFknJeiiWyGrsiRCV4WOZFgclyhUr+j/NCX5r0C3lE+
unBZdX4bkjfozDBgHCW68elzY+cPeLkwQl/QHVygw843+iLmOiVQGfBvnkbB2ns5ialYkxcxZESe
NLOph2fF4ohCPS14V/YDML0Z3Fp/0LwoB39PeWX3O+j1iScRwC5kAa89zhPlmn+dojQg9l3qjfOU
6na5aVeLd+AFlwBYyUaf1eknpdma1gfLaIj9Q1do3wwrODEN8T1efuRrvtgaGXZ81cI/kjYUo+rz
hgdJqtcYRF8ToXk+ibnQYbqrbDjzp4icxPRx6mqDcqcAVaPvLqiMLyLkijFV81LR9mjIenCw3xJu
+dJJQDZITykMKtiJYX/MwwYOaiK+qt0mFynw4Yq8wQbZR9WVlz/GDjamx1wtyPH38V9NRVWNqvtT
EQsMuSjWccti+SbXkfdON9oiJY30N3fR0eRfidsnwm7wQS3ig8wkcALbN99vdOHLHnoIJf//+pbX
DHsVJNjM9yhYYCSF+4qh+D+eMY6wc6VhSN3eaXOPcrt6yEAEwvJ2ulwh7mFqwgWvRyEUNEEACGWI
gI8Xwmim0GaLDFd75xK44zxbcuc8/Pzm73I7ibnX5GU5eK/xO2V11Yup+5U27nlXQCjg1aNgjYMD
makTBiRjLug6h+kMgBsbWTL8w0aZbKBmn8MCYMiDLXrrvCv/b3P6fLeu8SF7nLgSkONzsKROdeiL
59BB52sRBb0qGxsecRA+EK7XBvpJYB9lRKyHJRfV8aH8Z0hzJJBC1GsXZafdO8726hgeK2iM+CXu
/VUJXady68ZCfIKnQwL8oh579j7H2NYrxJ1uSj1GdoqN/lZIntCFtmy+FWXv6UetDOt9iGKKJeZC
e7+R86QWDhI//6AKqMdtYcTyG+biHwUjcZRjLY/G/QpH/mu7dtu8lASTvSO2kPaVr81XKPy+q8V/
cn1PQG+MppE/2YSe1uyQEpVT8keMs4FfvLQoQdGgLkNI9g/CIMPeqL1Yna8sa3tpWy3+tegxwaDn
RAZGq9Igg8NfyWewaA8E6F56bjYAIuZ9FYW8W5d7G8yHtaOeHS/AEExcAo34bm55+mZIWwKWK/Vd
HxwhJ5QmvwMtAR1dfa1h+5pCH0karSi4+rslIBcAT6PPCGKwMtEPkqq1SGGe+08LIPBFXEdkxVAn
GzxiXq5oG2KFrwGlgRBlHNQ8cV65wJyXUAc25Hube8brZLvObe8EOYgCEIjZJ3mKre0DQXjtwzEd
H3+MAbhM2WwTk9/9fTET58caWFStqA+fANCjwDTm5urf2nL60gE6RQftWQA5hn0T+0QuAbTtCv6O
W43JPDnXhEtJ1x9EeEAZcQkUtY8s4It/kHgjjRGS63GUmX5X5K0aQ2fOBz6S362vBFiaTMWS2Bty
cxxVdT+vAikkZMyNMm/luup4957XBBef6mwEd6nPLdTAYK9ZQrK6SOb5yPMdjnSKUvfz73OthNlH
JBEAtcpTAy3kJ4Y77Gkdqy0SoRhmgYTHGHctxxAzC72qnysKOOgBW+UDlKyvrFGQBq7ASH2L4arE
mhRrI8jjlmz2EFmjahwo767pwU7Ra5IPviJSO/i7i3dQdUr67dTP40jmMYKGsIqqPi6Q+SLoqqI0
hfab7Cijg4NY9VqY5DP1OnrVanHYht/BBkUdYhJF4sUW3cEem61hlFLdbLOt13U0qoBScyacXZaA
izDStStse2ekZK54lrF2u7t2VuNoQVbF+jOxueyR/vm5z7lfdJXwV5vWZZ6vv0vO7g8SD8QD9dgL
dhpD6zuLOwm6QxVuJedtlTzxP51+feYilFfkQlsVw/pJNEJ0vzUebBKhnyzE08aXd+4z0kZeeF7l
I7FjkRUO2fsFDme/iZ19UW7ZnXCdMM7mjlsxx8OA8SSfDxJSkqJx57sAri39eBtrszqdYvPkr/Yj
ywwRaWrhUEvxlMMtrpZF5JKp80JHKvBAgDRJg4h8Pi8ccx8B2gJ+wiBp3yCs+YrG3i/EYqCQJ6rx
n6QMAERDby1vTBmPPvK7LGBhkO5qS12fDc6dU82qVodoY5W7WXjE37XTN9xlCa/tHTSMEGlJpJYC
Go6BedvDfLpF6Pn6mXlSvAelWBKWVqDYYegZbbV2GSIzYfBS43luMZ0P8lAZiVWYjT86CuK6R4qJ
2/eyoNJHt3fUYLNBMNRGVl2R0PdM907FTtgbeSzIc1AElHQis5OP88P0gEwhkJVKs1PzPguOEhgT
jekWgbBTAZpQMoeSpP9kIz8NB1B2rtzLOSG9o8ospmWt3cnWxsBULriwMAhww4ylKq8e7nDTgrzE
P3No5F+wZo4O6qCk/uyIFsC5kmrwfwoMtfWffDbvASfMEIDsBO5tvOVVmQRvoOSRSFxlv8Teqacv
noe3OW7wcZ5z0DjgGFUnLwDLIIk9G2jGoWLygOrvN3EDT7WSdgDsz08bJfq/+rbk9v6HpokFMcEs
b8weh7rJUJe1H1x0BtWrvkDeVJ5eRAEx9kSzsuyZ4w0z0t93zb75kqDxuwR10+nhhho3E5MGIYgB
gRAZUTGl/tqPEAsA9LAD/oX9qwY0Wcz96X1tcFr8wDYVf/iFGMkZlf4oEqipv6CP1Tq6Vy6fdGVv
HbY3zCsvk6EcPa/5noB6IVX9ffuF+730gAfy491YCuvGlD97vfXxukBwfu7M0+LI3FTYK1/3GBjs
XjnpM0rxmNVTryBvsx6o0GF4EbhRg1YMX3jqBPqqYmNbQRNDxAa+89RXitOuCeDEOWQ0zLGqNV0I
iKZEakfvgWR89ubehz3sGH39kxCi9pSNsij5YGoJHJMcLf+8NBt1Pj9de0CUVxt0wmq10MWPoj3T
IczR6x2s63TbTAes+62sV+sFyrLLmZph7DoQfaahsNYKp7mfw1TTJnp0EvU5x450xtuJnZVAjzY2
5GXM809gVBQ6BpLO+WhonRq2RdrAMMhlD9MM1yNGjZwkezAGRRAxjYk8iuVRBxKC6lXcSP4TJt4O
5z+YG0wzLorS9UEPG+8583Qy4mj4InzQV31Cz7P7UMzcv2GhdqO6tC7Mk5EOkHG4dLbTHIOGVeFB
PoyPUOvgVIXwV5V7yeC88nZQSfTwsOstC1TyRsPFXqMdOkzj/CF55tGDiWQzXmBczO2e113G8xec
QB1fTEQzOugHFw3ORU5fDAB1fVOeyydO8ghKMxYDXSZn3Tt/g/HZuuMmDIRVjaWzHQC3xPV+wghB
PJp8owd3L0Ap2h8wjiN21gefQqDJoB7qNPQtRauzsPwOH/5SmLWCBjO6smqHwI6GaQFKZTA8F9wa
bTZJBgKCYcf2sxLFgHwO/to3yEJyS6iHjlFdXriCqJSwuza9wGWWrOs8EPpGTgdBSdf4zPZrKhzW
JikswfOTvUUdY/hTiWl9GtFbH8wjDsZTPuy1zSjFQ4SClONuoGDkteh4LcGqpnyEzucC3kAMIb4J
1cqmkIzrtU4BQt9qoHAUAeTKzy9tq0SqAClnE79F9gi54/TZr5MBmQmhKduGc10MtFwDnJPbMZsf
363l65jOjKES+x69k0ZnviBGeS5GUy++DsqJiTwf2ZB0olEs1MBn+ooRGwOGKUwMAsqoa0Q+Kv8I
0t8/cq4VY5cb8C5sdGI745IIVPyfbd7wnouCxfC+8zrbYXpwuO4tPrRse5xecj2qqALgsGYBz4Yu
4SojHIVN+xT4r6Lw2yReaFpT4gevAd7Xg3g8RyOj1Eqg3dzQ+0N7L57nV+OrRYCadVLcphGo7QSK
qiyHSuaQj50Rdm6iGOetdL/CzFJPbKWVPI71ueVHAp7sCxUv75WfAex/As+sB+PRjBO25Qixq+s4
lXLcRA7Y/E5qHZ8U4MvhUlQFRJUBEfbUsX3M/a/blTuVoFxDnoF1Dz0eys5q8skYxAJeX5GVT96l
gAVZXV8DztpPY8PfuGfheDvXcI+j/MraEvwJfGyzwk+Cotpnp6QDUDRTZFx9aYYhXg2J/3XnA3Xg
TJ+h9s4+9E0IwnXr60x5n11mU1Y18yyWDX9AkHypw9L09NY9fMLSgW/5449uzYNDZ2G9qE5rf2zP
bueJPZ+bKdsMnyJ/Ea1A7ikUj4JNTKy3AiDCvDpOMPxKQQCmrf1mWssyyQkDDioCGcMdcVtvaZyl
Qcji/+PWm9nZcL+FMF5XA4uHBO6sM/zn4nH1CFE8DXFuNbtpRvgeBaLjGp97ONS7WhoaNymV7fmM
hNncDzhiIhy9r58cd1XYNl6A39W3OMFJVVP/m7CHfJKRLihMuYCpzDOL6cWg7RPRQIX4cVAGRhce
C41Hz082tuO/M3nizKdm6+qAODBtTRkCGa5sv6RN/7OzWy+eH49/8GK2VeEulLSzwAJdb9RJeuBh
UgkUAtUdaakl6N57iXyGX8QYFZLFiPqzMgemPBv+D4wej8eU4/Gv/oBdki0w/z/ULWcasPKLhDNF
ivQcxVvhYwyTUwSZxJjwQtblWlFEmbu5QNK1npHy2hrFJG0Uxrq9ryyukFP7Qq+QicjwTADX3sXy
O2SKsPcJb+ySe1rw2klbKIL28q4Yvl3WtXvosmIahV957tAlCUuPxUL2pkbHCgM3otnh1a37WqA3
CDuWHtnhcAwtuujUTfU1HkM+/8emXrnk1fYTmz7wUy8x1ucP5j1o7/lxwFKpbuQ3r2DRBdQYcjB8
Lz2MYCzsNeWzrbmpou25lpMgVF2pylpZxvVN14YzRDsjCUoTkbKQ/Fp6DTwIy4ZLc205gWevXrfi
LfjYYzBiv++k4nxZsDfpGijSKl51h2UHe5+Q+wrjrVgJrBzxaZvSl16Pu1fIQve691AZr3XmRiMg
XeOsf6npMVzrauhYK/Wcc9tN27jkHE5u9mxKr0upMxspJOELoihg8pbp7aO8Edueb9ClMvSPMp3I
ppH5SubM80rf/ihnu8iGzjAQFK6P7/SYKeCKcCpCFIRrO5TtHGfIrffD+I11sG9k6AwtQFizBIvq
RqKtyoahDLeXM48YYAlpBb0P/0Cj7l5aoz9fAjekGhyjV1hO9j4hoDn1tVfndgJMrROy8qSjzVF3
Hcs9tRih5MJ6akswSZr2U7mt8eiA9bXLnVPQyASbdhWyLwOWqFITHjnGtmJ3HEAADNYDuM6xm/Nr
/yk5oK33jGrvDA9zByHmjnbI57iKCxkGw9LGyqidDbMu9RCfq2OEs2DI8Xs4lqOUpQU+wcV8nSSv
KgCVG4zm8URm+01POTZobkhy3rjIQFklLU7jCRn0ofeKEgejkXe45axQanBQoQqgbt53++P/hUNS
tC4JQ8MON0+OIdDEVtKplvamsNstXLMcau5mxR0B2sWf8u8e1pBpKlwcHuUjWOXVaaiFxQNwGwr8
o7jnASF6SkVYKaMqwsvRikhMNYq2z3Gblweqck9bsNV00VqGXz7At9fgW4pyZbVygz1+Zof8xDY5
XfAKnA0+BIg+0T7qGFd/KbQJQozrcihyQH2vpxaQFJTDkHn1MnWHWHM4/zfBHADFYjSTEb5p/Abf
JDraxAYrHEkf/eWa+2VjnAzt2QASKp6Y90gfJOOSdWZ7y4dIRKmZd/MYedfCoC1mAMzIIKHBqOD2
H6CDjsESytcMZHljwHSrZMPtYoKdDw4LoVSseBlNDLmfdHAMBi+CR3pozN1a8eUQzBA38FhtFYkm
bxaxxAiLxSYOiTMfUSi1Hft/SJk1nRAS2jB6mdl+HC6C+CXYLCUYbLHbmA19dJCrOJRYl5BOyBO1
qhXNb7SVCpwT9efrgZXy1ssWoPS2gzhcQ2DmmU0YXsQEZJEqUEh0QyjSvXWO040LzMYTIxfLb1fk
wRZ52NRqXNJdj6PXeBWpLNYtr+0hKd3yN04n5bT0k2ds5VIpfYBdY42P9gulmyeYROYzHxtk/eYy
x7jE+zh41Cu3hTlLhnGOL1joAAFhfIpYyfxjFWIezmm9YlLTHqDK+thm0soaJG4mQpOMmwad/7fJ
ld99uexpm+y9tR8FSKlR+DzKWPoVSV1IRb5yzVDV4kqzHBLYzYlgnxMZjs8PDos3l/daF/N2gnaT
I8p5BVssgSKThPbhWZWW5FdRv+1kb81M92X09YQDtDnTa4w8MA7J7rOYhKvaoiKZ1THwU/EeQzur
2daNQwm94XBnfLvV98Yw4nrgPtuZrCNCCJVug0yw36LiH3fZpDgKWufJgugaPOAO71WV0QgJnTVM
fzN+W9R5KdDUcMIZzH2Fi3is2wXgu77PAOAK0Gan1qu5mmgvF40vA4HbRagxo5nC5BZxXszUWE58
+exRPPMwHBBX4imJjWjgfvwvHloezAbSbblqXoQIsQysr/6KnnnERFXYDw3Vq6JLoDFLcBP67On9
1m5SZw==
`protect end_protected
