��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$R�蘧�rĦ����I��X1:���o�kܿ%^�Q���Ym�����n_|f`�h�I��.VW��Q�X&��	���a8k7�[��1�^�������T����x`�6�(���C��l9kUsA�"@�~��:6ߵ�y��
���e_:�f�2`Mp�6��m�ݗ�O^[COup��[�KvK��$=�QL*
7�߭ہH�)5K��	9?�\G�^�d+�^���H4O�cy�,�aS,& {Tj:��ݨG�Ǻ�쏈��/7�7ڄ_�� ϸ�~J�@�t�q=
χ��aW&��"((�'����p�j¾²S{c����Ͼ�$���;>�ؚ��f��P����A�:�4��f V�W_ނ��	�eu^2��S뎙>�h��t����b"�jK�+[�ɱ�н���E��EU ��LUf����]��_�^�x�"F<��lpj�mguR40}�6y{���؅��?h���<�}������0wJ>�{M��t`���p2f�9x?���,�F�է����D�a��A<�j�RPӃ����WL9$)}��7�?7®yK�"3S�d�<A�><-9���+p���[q$�W3c�b��-��$"��
mdT�|��9[T���1<gSu�o�dq�Bș���U�.G��A�Ì`;��h�4�٬N�FX�;�d�.�ƀP����'"�p��?����|=�FN�R����Yc*�w��{�c���Z~I�2�"##'����*�P�7��������:S�4���{U7�b��۞Q!��oӽ'��]�����h��Z�c��p�k�
�����������K���!�&�nFA���t0s�3b��Q\�|#1�R����X���D�������CY`�&�?�|���y��B�ݰ���`�����K�	����[���T7�4%��vlɄΌ&a��
(X4�n0�oՂ,�(��{%���d��!d���Q��D-��+�2��Z�l�CB����^��p�sa�w��
�0b�;j/�š���8�d`VԼÖw
�f%>l����UO�Қ9���}��K&J��؁?��G:�D��!t�U���&~�����ż��K!�/�t������JU�K��F�(ZJ����XY,�֥5&����h�Ρ[����PƮ��]���Y�x��&�Z�!���!�Q�	�L�%R��_�uY2Ql?Mq2��n)Ķ��W�,�v�X������@�O
�� :N�����l��s���;$.�W���>� }6	�K�	<k�z�V�鳻��lw��� oP�p�Z�G����BW�K$ĆJ�G��3��j��ư���׉4h˩�D��'��.K�t2<�����l�/O�N��퇚�NO���o~c�g�{-� ��6ݼ]�N�yg� �h ��>�]C�����#�<
g{�J��F�����r�캫&?��@z��L�zR9_5������t�F��X"e�Ln��]���m�P'�z���"[�����Ռ�m�bo��g�L��\̛)����	�T��I�՝���`y�@"Q=ޝ>c
f�P0�O��\�@Y�cD̓>aG�us������W³�䟛q1؅�yXC)�c��]��ը1��� ]��H$�I
����3���N6����K=Sf�d�`S�8oY���;w��g�o�v�m� �cC���(O�`������z $j�hj���"{b?�4F��f�I��➶��H�C�����;(>���f�D焗�J^OZE�h�F�z�c��7|^��z�7���cci�`�8�^B������Z�Z	�MQ�up88�}1���,�ĩ�1�~�0�5����0#X�=����V������x.�'�';��#)��[�dgg������R�D(kژI��u}/�ot�66�2�A������M��D�W�/XjJ(JZ�q�h�}���b���[L��񄏀Ƴ��PlDr��XC�7�n��}'_+���ɸ�x �~`�c��mef'��k���|����N�B��)�"����\���ؘʐy>�Yaᢸ�
Pi�3��Z�ؽ�<��H$�ؘ������63��=޲g�A|
C�g^��4�X����C z�s��2�����{�+��>�.��n�����:������i���(7�P���G�[�L&�KM�jy0��?�P��"��Za(��XG���y��蔙�Uh'_и�o����ZI1���h(��F�H�@._ ����d��Û=-?�#y�!�x��#�׆h���SJ�\�n����� ��,����6z>q:�!��9,��,nt�$��VMH[0�-bܺ�gNq������˅��ܤ����,R��^��q=�xD�����,Bv7τؙe�����X��G������R�h �����w��iY��O��W���\ ��Y'C���n�����)����&�n˳�pVp3��=�]��ĒE���]-���:O*cV߾�/���0����x߬s����9�(�!�䝁�͟��0	�9�B�7]��$��>T�Y�Pr�^�a[�~����ez+���ڀ�z�憐����G����W@-�t�&Pz�
�T�̥��NPo ��E���h�D֪&�D�/3��%[����V�W��O��pE�,���N5�~X�y QZt��J��$�ϊ���c�����U���]�%�(�v�khPeԪ�ǨNW�"=M�������iF�b`e��6���ʁN�r�I�*&�83��*���^L	*�J���r93�4}����c}�)ӯ}�m����|�W,�WcN������a^w��3�	v�Y��a:���G������p�<Rp�xeZ����*Zs�ft㻣T�-��������ͥ�җ�l��?ƚ�0�����ѥb�l@���z$�}�wF����P ���2 /������8�'��׼[�E�;�ԒK�D��d�\d�U��n�qP�ɋ)��y�a���V�AZ�� e Kz[��$R��:�q���[x�xߥ�j;~C����7c�R��gΕ	�p�ʮ �]X1��%h���!�~�ZU�ӄ��yVr�N�m��N|tS�K�/`����>ȿ�EO�b+�ʶ��\�c b����M2�����v�N_�}?��W���ܰn��x��<L/B��A(I�I�����CDF~r��pdg�~NkԲ�KUs�a�&1/&��<�Bd
u��-��q+��L�X;`�R��=�M��'�\�1�߼.}3,`Ĭ����<?W.a4u�Kފ+���U+{�������~��]��`��ǝ2}[9�X ����a��$��}�F(�{��L�TT���ɞ
h(�9t@�h!�/������HG��B�]a^L����Շ&ԫߘ`D9��0;��L�Q�u�>sҥ�^������8V�R�6~O�㮞t����f6�Ӳۈ�,�"�նi��-�EO��Z%�2.�JB6c�8Q�r��j,\d�i�ӈȁ���GC��>��!P��Ψ�!L��/��d�eƍ9>����f!��2x��y6�<���q[�yAy��`j��޵���:�:��W�}�p{�ih88l�	˄�frrP*�\.�qc��Q��џ�%M;�K��� 'xɝq�
Uw$E0��w4@+�ڙ���h-�)�b��1r�V4��r^N�-���M{��n�'%I�@*��s��|V"�����7-���3s�L����k��KlQ��ȊeB/�8�FP�˼ꙟ�Q�^�A�y��US0M�`���*7{ۙ���py�<�ִ0�_'�bﾴ`�*<|��יj�+{�2��Hy� ��\+_@g?�<��(iG�j~5�_Bm��aL�����������G�H諟Yߎ{���1;_Bc��˞-�l��U v��a� ����r�xi��������| @���
�N,�k�:�c�O]�y�f�:v��1���1$�j�Q�V]e��S�,�%ݩ����!�����g�S����:���gz�)k٘��(�{k �����H ~�?����vo�G}�(�k��-*�s)e��-���X�Ϙ]:x(��d+�7h�P|w�zo^��K�R��b0�3+4���<�Q���A�`[K~jz��u�V5�xGeH}^h��((�	�z�T��O��9@�y<���P
E�S��y`�Lz�}�xeQ#cj>���A_�[#Ͷ�3�HP��/�r�:��R�~�� oD���	N�E�ŊR2z����sNz�}�Z��3���Y�į�b�E�����iG���ec�s�÷�eB�H��u��he����ihgLYIi_n��$�M�2�8���������j>v�u	ߧ��E��г�Ʌ�P:�2���o�����2���S������%@:=pۀ6�{�?\�6�g���ŷUɔu�w*�ą�l�L��豫���U:�;a�>�3�J��g�mO3��\�`�谬�c�Y�S��w�P14����J�%ҩG��2�l^���)#�� ��)6�>(D^0�%�|f���F�iE�J���^����BT(��J�N�nΫ�<Y��%�D�z�� ~+��vX�T��E�Ƙ�:�=N�~�DfK�Si�����!
^�Ь�Ѿ#�{ߞv�Ԃ8pe��0���޲��L%�?��nd�竳�n�2�I��F�V�G��Gc,��C�9��=��ªb!ؓKs����[x�7r���e)�y�vb̰6��} ��צ�i������D�h=�K�A�aB�3�ʭ"x�w��=�e�WhaPy��,�ɑk������c2�7�-���%�����/����5뎥C�,E�f���a�`�Nމ�Ph��!;3����>0�@ �%D �s�q�1�6������a	�ծ!�!�+#�^*���Q�B�����k��zM]�@�h9�M:D�8��@�����tJUZ���`�	���n��.��8�����Q�Խ��؏���P#螔� 8,?+��ec)��L_���p�������F��
?,%�aܟ�W���+x�]'��������O�p��
0��s���|!�[0
o��"֢f�����|�\Y�&�m�!d��3�⣃,�9�<ğ;�ٺ�ĥ�1P=�s�w�XV�wV\e]�P\����a@��q�(*�TC�6騖E�;��wv��|P͔�M�eM\L�&		gx�挬���\��:&���}u�i'�X��/i)�x�u�����H��G�`6��o�^l����9o��n���CTe��bdM����x ����<՛���"��W �w^ӌt����%�+6�������Y��c��A�A��S�E|i����-U%�g9�_l߈81�'O ���[��| ���:�<��u�f_5�[�3y듁�É$6w4���S/u�ZI����?�{�j�| �[�l���&��We6o�;�ً6-pJ~|��?�X�N�(�����c�)�1o�&��,�il���Y-oǖ�i�A�Kxy�7�s���JJ���� fҫ�[��35�L$`�wn:Ml��>4#$�հ]<���L�ޜ�uT��5rOd�|�K��QO �#i�AE=�&h����Z�f0��2��5�z���b�*��v�| �g��o�B? �U���0=CX$
#]����}���ÑXz@�]�_-���U�b�a-`e���1j�W��ǍBs|&o�Sh}�y{�o�Y��so��^�����@!�u��E�}��b*.�P�"oi��]��4�BB���z3��+^����
n�JG�lV�)��ZT0�>��mo�W7̪1��V��a�g>����m��I8,h��L���9�{�q�����G���<��M�mj�5�*�@~	%���߮�ձp���$�W��N�P�a���vu�ܴa^��� a��I����ms��u
��F ����}dʿ�� ������1U�''��n"ac٭�.,{Ϻ�[
�nxJ[,����%
{)���㹔�����-�熒O¿�T�xJ�PP�M�_@EMT��K�����*��_�j?v ��-R��7��WjE�3���`�G����{{%��/
^�E?�vC�������p�����4K͏��gŬ��?����� �=��qM��'���|_EV��%8"�F,�u�ڡ;�m�t}��mo��+9*�M�`�$��B�����ߋ�N�����xH���DB�Z��NnLl��� 뚵���Q��	������S��U���������U�\8�4�>�F��!ihR��c�Y�͂ZV=,���spS.�O�E��BBa'�R��?J�������~��y^%��h�6()
*V��0۝��04�Y�ZB��h�MX�����7c:�Ѹ�q"]�dC��}�m���t��;
33��t�r�0�N�0=������,L�����΃�nx����-��R�$��9��0uƞHOqX����Y�9��&Ƞ�|�@p��CU�ˆᚹ�wA\ޮ�Q��1 �j�Ĵ���	�:O�$��
��w;ؤ�c�������Ѝ�SU�  ��m�t���t�]K)cЮ3�V�ذi7�1�.���>���y�����\�kc�˔k�U��׿W��P��������,�.�x�:����y�!G2uG�V�*���
f�!v��' �b�g��
4	B�jM�Bn����z�w�V}���2�4o3E�u�弟T�$-{��= �!�]�������d�DɿB'z)�L�B�4��Ez����jʾ=�-��V׸XYī�t��2�i9����)���[�� �Ч���'	��+�g���o4��cIy��������Wz`������6�U��>�r��-���:��d�Z>qJ"�':30A½�����C�d]�mi}HDk[��S���P���Lm�c���l���6〘Wlt8�59(LR܎Z�\�fg���/�,'F�C�9��N#�b�h�Y/1 +V��i����A�����3`6��Uhw�.�t_U�;�eA]�Y�4^�Ľ �s�<���ֺ�ũV��uͷ�?��&J�6�[�/pq075�?�-��{&�Q5< �B���t�T�X�\����aE����?[d�靵�E�n'�}� �^ F6��*�P����
?�\R�B��
U`*7�[^��K����nHxO�UQ��ō�Yh,����_ �,p?�H����6QԠ���!���8��H~��|Ne�]�s�o�i��?��K�;��NY�M����Q�:��\��c�J�����>��
�xKo7��:����UF� �4��(t��~�Uk�ä���:Cn�[5կ(`�1Ш�B�����=)Z6{��wǭ�`M*�Er�C�mp�!-V��yh�<虷u_D8Z�v�;������H�Z1��	w��_6�\����z��g�Z�U���o���c�R�F�C��J�{W�,懽��L 
P��)�?	�'�&=��­���y:,��I�����.���#�=��|^���6����D��z/?���S�e_�De���[u�Yى�TQ�7Q�J�}h'��U���7��������'��:����O>�3*%��h�d�ֹ�m�>%�>R
9>��(�Bt"8 $���¡�����5n'�����׸x�ł��tϚ) ���4=Ƅ����P�h�l�&�~��V�#�.N��z��[�'8���Sm���MQd:>e�͡���Q� ���~�ZS�Zt���u�L}/xñ��j�2�#�y\�h���<�=D���Z�����k;[f�9PKΡŉrW�k.[T���p},E���>-�#��"Pwt��4`צ'���^�h��*)��~�W�;�o(rq����7�z%���`p��%�v�L��+����P��v�!�ԸYn�� ��M��![�ON�rH��	��'5}ݢ���N����5(�3�T/Tc��'��Y�'�ϣ(�<�d�bqa��'g�Q��(��� \��Z�oOZ`�+��fD��b�T�a>�,�^�9���ԉ�C]�-y%��K�*�(�[S�F�����L�u��5ZA�M �f�~� �������=�0\#3�nb`P�Řܽ��*~�:T"{�hHq%GS�O��) �{��2����ṙh�&D-�?1>lz"as�_�1*n2��R�l��R�����6i
�J���K���� hc�e��k�N֩.Co`�Q�+8�ř)�Ac_�O=��XL�%�2k�H�%��j�b�j�=Ѱ-\Ղ�u+��ȭ$���t�r;V[��/�ź������''�f�"-\R��a��+�{��g�Ӽ(l�`���L��c�̠����,�_��`��Au�o�XP�?aU�*�$�|�{��l���ׅ'm[�h]g��gK�4{`�+SO�eL�_(�w�;���wma�2Ks�����{zv�2ntӮ�rG�\!#H��ԣ��F�S/�Y4*��ju�N�d\OJ+t�<�����b������;�Bu�=IG�t�[�Q(��P�<�3�{�}A��Ϙ?��5y֘�&���%Ҫ<�M^��S�����K�{Vb�-{��|�����j�bq�E$����Ta�r�+o���L����'��X�5��>�PYWi�I�#B�J*���P���R<����J�<8�,'�$���_�cj�Gʄ��v^M�/z�"�5/��hQϊ+�ޯc����ǚS�,�Hj-��#	`���q8�?�~*\7܄�ɼ�.�{�	G56�h�ٯ�R��p%�o�hfңk������R�@�Z6"C:r�& �{r H�}	�����#HQ����}:�_�䣖�f�*N)�Δ"�GL}�|��K���tt��?�-����A��w�s��٣��򸐏��#�M1�K���q�����3>ʭ��Ϥ�:ew���bA���A�>�tCмږ���֨2'>�bC��+\"A<tJP?&2W�G���o�¹�����O��z�d��pɇ���`J�|�J٫/8�������!a0��!�^���Z�(����<y��R�^~9L�PEJZ���j���j�0����wM͐,P��b��ƻ"D�3.z{h�-��p���&�X�|�#�15z���>L�þ/��M3atS}L:�#%�c]�א���p�LL�i_�����[�$TJ�W��V�3~o5)��c��3��M�3��b@���be�.����s~x���>)���fP�^�&���5�OGzE�� ~���D�F��($'�����i�����,�s���/�xQ7��'U�WF�>�\:��+�Y�̗0�
&м:��v�9�x	���T)°�d]FHQ]Ěr��?�Y+�ۍЯ}�@�2�F�գ�����:�+�B)��G"�F<!1.��kLU+ 0A��DV}5�=y7�d�_��r6�%v4���2�V�	�H ��& %��$P�/	�T&�Ҙ��Cdd�oz�Dnl�[(������V�$6t!�5��/"S榙[�2]��
K �Y�����,��^�������{lO����߶�\�eH�~%}+����=	��F<��+��A̤P�w�^��N5{U8Y�OŠ���r���ѻ���R$��Z�xZId��~w=tl\��Ƚ��8��b�|p����S�ܝ�=C(�!�4�N�����E���f
�I��R;� ��>��:���'i��,w"��`nAGݧٶ����y]�#����k�W9a�N�#��-���˥������C�j�#�z���1�L��g15.:�7!<��xj�O��h�?a^G�����|�b�@8�W��
��'��L�xU2�����5T� �b�xG��k����m���x)ŧ0T�T��R�%!3�'&���?s�]�Z��
��4%	IL�Dpb��jE!�i.0n㟥��n;yOă�m)5cvu�0{�
4�NFVܚͽdO�\��]���띵Pbx�\�ٯ5`}C�;�C�쒙̓�9�"���BcyH��i7xd���'H�ax�L�
 �U�mSJ�Đ�Y�|���tj��'q�#Ͼ �CyTtl���`0�5��C�s��q߹�f��\�謔h�]��D�:���{��e��&0X�>i��Ɯ���|W�M[�����R�G2{��p�� w��� ~��o��d�(iT��f�q����
Ao�L���ϣ��&"�?G�T��b���Iw�#���Ky6	�_u�>o�u���Yp���W˨X]�ԣ{�pR�	l��cɺL��+y�'"��Lx�Tj$���v1��|e-w�.u��pyT}����8�ȼ��R��Wh��F�(`�n��z�a�V�����0*I�e��5 L������,W�p��.�xc���S�F���׾����:�"9��NZ�x��+���y~��υjL�I.\gP�.�L3~�0*���ɃۈמM��)]c�g��Vi�4�
$�~a!>���#w~��C��ɞ	ڠ��6�H�大~���qB �ĄΘ����Ǜ3d��I
����6����>�Q�
VY�^Ky),�9|�6���6�Yㄋ����r�w?]�cQ�{L����~�&^�?C���R�Bh��xp`��,\�?��YU�3m�K�(�A�VrN�([���˨��Xx��szK���b��@��R^��r��eFCC?<[�l8:�~C��h�S5���&�D�5����Q�j+��	��Y�����ߡ��[@�M�p��@�O�rc�E�Q��༷�f�ZÜؠ8�n��w;ri�#�2R�@����Y�0���L¨X7�µ�--3
�w{a
=܂Y�L�T8j���R�2 ?� �_��0��f�u"$�g��?��
?dîӪ��Mi�}Q&jF���>`T<)��5lU�}X�[:,u�;����tT���U�BX/j��G
$���s;�l��I5JJ��R�'�A���ǝ�z�/DQ}x6H+W���RC�Q�Ϙ0�`�@N�aC��"�	����">A}H�Y�����St�:�ό�X�U��wK��65(��`�9^L+ʔ��׿�Yer�1*��ql��qq]g��ƴW�����ؠ#������2��rR��ܸ�v���ex�V���L02J	Z�y���-8%Y3�
�����J�K�s���O&�ؕ
���71��Ƹ.߶�� �3Zإ��i����X�3�S�p�hǗnt%R�ǱYS���7�Z���IjK���r.��M��7�c<mI�9-ݿ~�!l���
�x�\f6��O�s��)�v��WT��&r�)=�A����-8Ъwjv��ױMho5	�6lg��C����`1:��R�Dze�a����ir
�WS�Z��HXq��E��P12Ea��Gv]�W'��@�f�����T�������������B�d�qߊ�k6O<(��n�3�sb���F�nq��]�c\�:�>��o��cXZO�\P�zD$��'C<��l�,��!�yY�ը_��x����S"E��ٙ_O$#��T�
YJ����@����ŷm��	�M;5̀��@\���+�cg(����IrЭl22ҙ\�̎5�'O�k���Bsg�r{��De?��``C���8�\R����*P=Zd<���;����Cۊ+`&R�9��7C�3d���zS֡��Q����o\�M�H�>"Ͱ/��pM�߀�uh7�a��k1�/{wMF� zNcE���\=��^�nMC�oZ��=�R�i�;���dm�וQ|w\��ȓ�����%�����=��s�*͜
	jq�NCq�]��������"�rBE� ����P�2G����V��y�����k�F��=e�ڢ��<��O�'(�8.��b�	�1�����-Q=o��J����Y�Lh��۸a������J�{����l���/��e�#��хMs���G��`7����;�������9'��w��۹��vu����(�/LA�|��Y�^D�?"�C�2x�J[�XE��_b��~t�Pa|P��~�ލM-]��~�ƷM��E�s��%ly+�1Wt`�l��+rs�1z���,�5�l>�(��l��
������kVp��ԯ�8\j^�N�=�fo��Bv�n��_�{��5.�5��|�ؿuP�"'=͡䳒����}��e���G���A�-�n��m����c;�Hܓڿ�4J��O����A��d.(+��o��y}cی�Œ琖�7���B�6]�D��0����D�P*��7�CCG�8�����*�>�o&z��`�E�\�Ө�t�\�~�w{���Z&RX�/��9�����2����}D�+M,-j�.a�ZP�!{Tv���e�!��+�����h�W�cN��'�e���r)N��t��ՏF#9�w�C�^�e7�_oH&"�7��k*��a���N��i��D;�,c��.��,�ֵ�R<ZK;<٥L�Z�j��R�_l�y�6��S���<�L��#/�М��<�R&Żz���@� :v)C�H����b����9T	L1k���ٌ����"����T������ϳ������߇a��G�k��m��w�a����,�[��_��IQ�"5�p�^��4'��+��n
X˲�o��h�l΍"0�~��d��[Пx������RB�[����&T<5�갦[�l%
ڞ+�Fes�pc���=G#�0����W����2�h��>��fa����J�"�}��`�껳��Do�D�AݓC���،`���^���������1(��bW�+�ĝ�+�#�������`��O��Z�P�9���R�6�\�#3q{CO,��=X�`YJ"�'� I����T��R��/>EP7��Th�7}�u[�g��6��&x�?H;�]<�R~�Tޡ��z�=�dq�@������&"�]���l�s���z�UUj\F���N����F%e�E��f�^ֶ��-��Ƀ���t�7>N�'=��;�a]��x����>���!�o��׌����ɮ� qY/qD��}#�%�d#�f60�ԉ�'��pxa�N��t�u~zX1�H�,�|~$^�>!�ހ�E0M#j�u���Eq�\3�)��Ge�4`��[�o�(�%3׋�H������B��:���h:��@��f0[:�sX����@��өp���^��IL�0�S�2�A���?
��m.K�����'9F�A>�(^r[�8d���l�-`mh�������Rq�&�	'�O���H$�,���!�*9z���@��#iti�	���H���?5�d[��;�&k���hx!@��������!����$6������/`ܳ�x�4:�dx��Y��8�X	��'��[䨉� �L��jp��	���q�A4-	��{$��l��w�eu�1�q��
v���B�꽪W��D����[�b���1"�T#��̈Znr��A5�����"�r��\7���c���F�� x?u�h�a_/��Z�����"�	vh���B=k��o�[Ǌv��u�5���eh_��甸68�� b{H�:Z�f]9@8Nf��&�ȿG�U�1ک�ܲP�f�ߥ� ��+1���y�Ԫ	�<�P�a� ��9��X`�ݺ�ST�b7� �
��p *%�:CH1�ɚx�V,"�0�ԫ���h�+��y�v��P���9e�?!�xg$s��J����w��:_�4W8V� two���se������g!��\-7d0�~�!e��$X���o$��E12�I �ϭ��ʕ�XC~6�7X5��Aj��*���B����cD���[$Qj�HGa��Y�eHS���L���+2ݬ�6��5J`�_�{q��y�o�z��{l�k,p�~�]Ӫ=���H�$u�nDj45�!3�Uo�<e)"\#�j=ƺ�Q�S\��mz���"���,�����}.��!q����B�*%��|�T�?Ŝ-~c�����bz�3Ȫ֖l�������_3���"y��y��g�x3GTկ{P�M�K���D�H*�O�]�B�t �F����=b�NYJ�g"$�F$+�K���\�'\�m�G���b6�$��m���^����)�5��6��"��A����oj����_�O�v��b�euT�,Vrx23��ё?.G��$|u��~��%t�&Ug]��H�x�y�l$J��;!�Uɓ���&�B��5�/�&��#� J�����؛��do�5)̟;'��zt$��/)�M�w�꿷:��C��;C#������NQ��|��r�&d�%#�Y�\N+Ԧ:�K��=��D���;���p��=8��� Gĭ�_/�_cT��*BE�r,ȝ���"C΍^w��O�c�=���ڻ�		��ne����ff��^m[iH�ra�"ɍ��/ ��f�g�O��iQΊy��#�?��G��<]���fkr�k�i����e�\G*����h�!%��z�1�"����)!����'���v��?��L�s)Ѫ.���$h�Q���^Gq�ƑnnD�_{kw��O�9�;�H�g��֙F��(	�˙U�4_.l<�!4/�A�{�;�Y��Y*����(�SmD�шl |��^ƥ$��c��"?�%�H��?'_uK�O߄�5�����D�mv�2�w���O-㧣ri�@v}���ɽl0�;���>����G/�R���X�b�9L&h8\e�S�S�O��;�j��E,٫Y�vDj��|�(���?,Cq�z:]�P6:��̩In��w6���	���(�i��&��F#g�>���Ŀ��TK���p��B-{��5�"�}5Nr?WCV��5�Z�з��T������S:TW�D1k��c���r���v��Y��{��a29��S���8ԙm������5���?�gpV3�j�������j������9͊��4�߄;��op�m=���&^�����y�?r�Qͺ�	N���`[ϛ��ym^���$�p�����/t��QA��j����b��T���.mC"��R#��p~u�J8�����٩M�VL��#�>�(?#������}KQ�
��H��}�n�3@�(�[�������� p���Z�'Q�g��T�`����ھ1�8�u���&ų�,��Ɉ���xǢb���A8]�cthسIC����Yh���k��4+M9���^��-�L#(W؂�����hg��
,�^��Y]��w�Nw�I��^r$��>�:Zv�"�:��z�b�$9�&
�=ݸ�n��Y1U!�S��D`�ϵď``�c�ta�ى��]���s&�#�_��]=M:�ۺ8.G�]s��e�B����>E��)�7-��q�$�/���I�&�ฐ����x���� �똓V�����v��3 �T�7���,�;/���SF[4�S^�N.l�ƽ��`��d�\6W���x��ۗR7)�2��7{gX���(��	f����@5�\3�0�!5�)����.ٷ�]7�Yb�Pm�W�#$8	Ex-ђ0�q������Q�ҠKJg��+�b7�hN�����u.�SJ��6j#|�҉��ת8�<���d�E��t�S2�fճ�z�$3R�x����x�W�1��ۗY&��.�rVTS��ɰ:�w"���2#��m�P�A��Y��~D#�̺�48�(��̑�'��k������ޛ���׌��#�6t���<[���pt�ԇ��2tn�]�wV�n������<�Jߌ;�G��8p�׺�mj�,Z�?2�q�-�����}T��#�f
���H�ߜ��~�o\U!r�3v.S{����9E�"����we?_���]A"/W�%Y�2����VKa��4i*���L��c�v�#���-k{��5�(��N�bY���� ��lPأ��|3�ֳ�����A6��1#s�0���\ESX��vUe��o/�+V�c�F:����*4��L��T۾�z��Y0[�"iM�:OV�O�0}��mA�vҼ�N��'n��1-g&��t~O{˹�$o���T�o?�]`ز�5g"�eB�C���X��ޒp��G>xq��|����]��0�%'�}i���ΉU���ڛUΛ��*ƴ9U����R�����?g��9�8�飑�')~���w���uN�=N� �*�xu"G��i���#]�[V�*�>w\�4�w�Q!�R�DQ���Md	$�3Q�kZ�e�[���I�zMjL*͐b�(�Jl-cY<����F�3CC����'(��˟:t���Kkv�`ص�?�,�kҜ�1E���}i"H�",V쮼�T�Vc&�ͪV-�Rp�PiV~4>����q_W�����.�����L���>Tn�!�y/M��������B�7uY��/{ `_�E���OC�(��7��� ����a��7_�h�� ~�Xwc�x���et,x<��wx���|�(�!⒎(UՁ���E�V4e���������n~�[z�?������&���T�7��<˞�4����e`9�AB�F�����W�^��r��Q]�lVK�<��g�*�vn�c�3eq���،��NBM�P�UO��>2ΧY��i�p��B��Dy:��y��ќ�e��������B4��/�V��(o�����Qd�E<anu���sp�R�ј�<��2�1��w��5�+5��~l�~���a5,$��!$��5０�$����^<�Q(�5T0��K��l���ޭq ��U�GP�$U���zq��>��z�עx�t�H��}P���t��3�RS+�?���=�d�Nea�ǹ���MN�(����}����։��Hv}�f�9�?I�=�� �\Z�熥]p`v@א�䳞ϱ�a�S�7�����q���%x*�EU����Q����.�%�Y1\)�8yl�KڜÈ$_=9��j7�g*��M��wroA�h��2�[u��i%8c;�{*�GÏ����_�:�~\C�����e����`�F����7у-d ��#z2A�ih�A���*H�`Qas�ak��侾��ǅ�K�9b��l������M���XJ=C� -�4騨	0�c�<%�y$��F�r5�k!(����B��М�ji}�"B�UL ��c�kY*�� Dw��`U�n�M��aW�a���dmM{��t�ПW �x�`���ذԘcK�u�0\~�����;Y��e�t4��6��lB`��^.���������>�#�4��Z"���1��+��A��̮��U����u=��e?��\I�<\�Oe��Z+�I�g�-[:����B���Cb�lA��Ǽ-@O"��I?���^I��#+_�L�N��3Ru=^z��#`��=lb��u���'��@hn�ڊ�L��4n�˃7�C��!�Z����$ҙ��v�A0�^y�քZS��+��zҧ��	�r�<Ӥ5�zt%#�+�G[�<���b�-��T����0^��n���PM"�v|��ժi�*��!��r�W�G(��� e�E�`�g�A��J�إ��Hy�<@T5>3p�`���6�[;�����&L�}J��nNpvuB�� �g)tqx*Dm�����ڧ����{�DA�VN��ʻ!�C�YH���s�-�릴�%(�U�HD�b�Y#�B���z�1Nn8��
��I��Ù!�O���mr��ð�¤U-)�DfX� E��� �6�ѕ}����[�w\Q�m�<(����q'�$H��G)R<��I�% ��o��X�;����P�}��r寐5fŻ�:��Vx���?n�[���<|��i����V����� h	8�i���;�MnD^�#n8(��E��V�
!�b��;1P�W0E ��$��Y�l�<�*#K�UXGK���Bc���-�R��@� ���~��^�N�?L$篎��l������z8�w+�ŉ���&J5�>�mxr ���8z���v��z5�T��ȓY[}�S����_Eg���F�?��x
��LS"�R8�"��%R�q��=�	��bX����jAJ�<+F��3?ر�Ao��⨹���b5��f����ty���"|�..�Dj~�GӄE������u�cK��G1��=�:!|T�ƈ!�HE7io��|�n��gT{A��$�V��>�K���S��h�b�c)��OW\n���s6r��i.?��8��/�V)���n �{=rlIV������S���%�D� ���&p�ӊ8X�2f�6l�q�k�L��27�eK�8��
`�?v���nFx*��b&.O8)�ɇNPj�/%�w�_-·�,�7��R�֤4a>����.����L
l��x�F��&m��A�uG��e�?E�i?x�#�LX���ށ7���6�C\�m��Ǎ�P'M��q�%�["&�e���H����WG�h�/�8>;�� ~�
r�,��]� ����w�ۦ}(I��h?F 5��FV�ۈ7����h�\�V5���6�>�?���s���bv	���)�?��������K�5�n�3yj�q���:�%IP�1�&
���8�G�u�?�Z�Q���j`W���>ر"�9��j�:���|���#�!g�2{HY�5�K��;�ᄟ�`�(�A{���J�����p�0�Q��ׁ���I �G���#�hn�e�����nH�D��P��;��m �>��Η5S }�3�v��MK��3�Q.�@�)]8?�W#ș�ͨ���	Ed��h�l2/�nb~�0+�rF��J�\���_��h~�Wq���|����NJ!���V�hL��?P���%V&9\���B��e�6��Z������������܍p�>"���g����r� R�<4�/�����@�:���sl��g�0�:�=�H�Qe1/g8=�W�����9fB.)�8S\��Y�����8>eDp���#:��&b����8��	�0���