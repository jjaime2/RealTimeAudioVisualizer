��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊b]{s�`���G�W��' �B̦B��yE%~�����+,��4�#��s'�v��v�.\��]������JBL��2Yt!Zsk���-1�h8^>5�Z���DfTo1�W������^����E�_�x���;�Szo�6�L�h*�>�*M����o��O㛍4^��(a�Ӱ���B��a����[ 4Tv���φn��!Q@����b]Cݿ�%ot�"q߶��#��(��.�8��w�9��5��[���%^B�_��;EM#�E4��/�]$C5(<�vn�T�[����Dfu53Ń.O�,��<�,v�Ze�EdX���"L��dpz��w�=e#���sG��x�sh�Ē����EF��A����O�i���[8��y�z�T풼s�Jr��{�Vc�U��i��-��H
�y�`A�Cp�Sq= ѕ鯢���1E���z�v�L����'|��T<h�fQKm�c�l֕�f�w̏�b�2�s�iK�'��; ?��'<���Ղ\�͘P�3�q��uƙ~���QJJ�% ���==*$3��- \���j��'4�O�������� m5:��~2Mʌ�����sd����bk@Wf�Ȏ�f���%�C	N��o�����\c|��A�u\�H�wJI��� ����BcX?c���\v���o�ge7Z�,����%�����r�����OI�#>�ÆX�M_	��I��I�n�y����<e1�	35�p��q�D,Y���`Ϙ~�X3�I�-p�VrX3��`Z�� [�?�n� �쐅a��b���k�� @ ���*�C{4_�K�X���s�C�����`Fg>֢��c5}A!`O(�dr�<�������1�!�	c 7@l�a�R�����AA��?���ӵ�j�}��b��?fO�z=�@`x��L�u�?��h{��L>�2T��ڳ*��mx��В���X|F�ʄ-W�惰�E=�T�,�T��,���zw��->I��$'���hV�ўt�3��蘫����SiZ׼GJr��&꫹��d�X4�` �L����
&0sx|�c�v�_6N^e����k�Q���38���_�n�r����<����v�)����W�������T����u�XS=���YA��D�U ��c
"�L��4�����k�f ��k�G�ޕ	)mq,X���0��[�$�#�S��d���ɜ���[.շy��4k*1I���D�R�[W��n��q���s|PE�w`=c��'-�����Gh�GB��a�?����?�̤b��Ll��TQ�6��>_�Ls���<���
��d�O���G�ji��b;=)**s=Բh4��L���=
C�!�H+�w_�O�l4��!�P�G�%>�a�F��~g�ͣ�xUNi�,�λ���M�l����2l��0!Z�l�Ų�[sS��З��gP��~s��g��%���v�����M~0�g^嬥'�8b��Ʋ�{�g�υy�;N���4�B&���Yj�1g��>�}?м@0�c1i3��p�D��}<q�F�����������zw�g���<�����Ύ�ˇ���̿k�8W�:R���r���+Z{G�E�F_�p��pb�,^?���ϸ�z�v�i�?����e�C����E��!~�a{� �BHc؋ mۛw�2z/z#M%<�\Gȫ���f<Ͱ��+���	e7ʴ�����,8u�pA�/�j�h�P�S	�-�����>�|����;nf�f��߬Ỉ��U�2�6���
�p���*��m7,T��]�n���i��7�O�|�J�VZ�Sm���4?>Q�(�A�pjr�Pp��[�8W�R��VJ�L6i��ѵ1��A�M~���Ru���3��7 ��z)�wU\gnNI��(�4_>.Jҁ�ȫm��s�V
C���"��T�^��� �М��˚6Z�۝m\�-'w� ���Gw*ح�/�ӿ�x�S���n@*N�۞���U܉�/:��mLP*^��V0Ǝ�;h]xd7r�3����z	�v=����}U)gqǙ���ʪz��;(�ǭ��U��`���� �]C�a�D�4�(��K	�X�F@�r[�P�$D�����&��3�`��� �/�{�1�j�ګ;.��M�h��,�mn�����4�
����w#=�����.��l�GDWv^�M��b��P��lе	�O���P�ki| �E�C2�G��Sgn��=q�h(�x. ��v�B��=V��hQ3��;��*��2J�D�����z4��$"8�zt�6��&��;���Nm�������g[h�	x��Ã�&��H��K�S �f��Q�ѫS���2��`�O֌)��&�sҾj�e�% �@�Ǧ��}8Do�_�*���p�*�#������y��?
���|/���M���o��M�vPޏy_���8U49���o�|�D:��ӹ���L��R��5��D>Q42���M�����٫�2��> ,6�oz�&� ��:)R����r�,���!P&m�ݍ������p�c�<x�v����d��q�(��C��[�c-��~����i艨��j���Ǥ��G�t��U�CK���T��U�?�������Lc;���.��D+�v�:~.���e,�R bM:�I�1��һ����.M����YO�I�5"i��՛�߭���9V���,� �$�!p�VSᘠwt4$�iӤoT����F�����3>�6���Z�����_<k���&oJRx����)F�3�/<�ܾm�{g�!C�y�>��물5���H3�iߎ�.�/{��~U�i�"�Y�orN�M;>����v&z��7DM0�p��)DN������a�}�i �e[�y�ChGH�%�^���ϭŵ��x��Ȱٜ�>�y�$q�Jφ���;J�&"��sC�B�dR���<��/ς+���P�����=��ڍy���O��|d�x�/y��B��Lt�,��A�s$��!�)?�"��no�p����,��@sZ@#[�os�"k<q��0�e1^�^��k��E�K�(�j?hȧ���7<���nZ�Y�P�5��H�-^��O���>�R(P&�=�1.�,)�R�����t���N9hg^�l�O�P����v��.���)|����M'Ai
e>$��a��bE�k��͔�*�B
`�{��?&߰��5e}D��1�[�ټymQ�C�NckK]��RO���V'"�������]��=�� ���g�(��}���|��A	��ؗ��sˌ;0-�w�����rԙ��'�O�����[Є�2���+7g� �<%��B ���� AiXA�+쟋I���`3���7� �0��VQ�LO�}�"��!���d:��GްAz��'��������3Ő�&�0��+�b���8��:^Bhx&
�R��[��a���m���Syj�F����+�V��l���B����5�x|2w�]R,��"��j��Z����j�/o�0Z"i��G�c�3�uoD�e�xw|�v����ԏ��ƫ>؝��<�Z%	��]^��HZ���ӱ���r��p{��v���j��V�N2;#[�s�뵲�f7ȳ!��Q�;�<auOB��.��^k���E7h\�c��#�Q~X)K�F�{u�!�]�q�d����_�>��Tu��STc��$��^M�@�]��>f>�g�(4����`�z��ϴ�'DJ+��
�P���߁E�
������	��5��� x2V���0��i��*4O�Z@�����`;\fuvE�	��X���z�̰�̛��l���f/G�JȨ�b�L@��V���[�����N�E��$]"긼?h�����~{��D�ÿH*�xU�CW� ��;|���	U�OYV���Ɣk�B�Q�öiSzӽ�yUcf� ���M& G�7�|,�`W�����7�(�
È7+�<��ZN��P{_�k�m�uq����n�,�q�[f�<'�E6�'��ˆ���S�./�s�Dy����W�ؼ��BJQA������±�U�L19q��;���v8��V�A��g�f�#4�ٙUd�q�PJo��J�Ei�V�2{��1�%
ݜ���w�X� m|;����e���,��B�Q��^ٞ��C�Dx8��6�/��_��DUE��\����SB�Ұ6}i �Q(x�Uq���|�KQ���عւ�H�"u��1���(h�?@1�8U[X�������[p���t���D#���:�.�{[,Q�} ���57��"���[� �����<���F&��R���0ܭ�Kg��UJu*��M���L#�Q�Y+�s�q.��Κ �e���ѽ)��Ȉ��Ρ�y.p���jĖP�*�yFc辧����B�0�]�#�ًt��"6�Ɠ����u�w�1�Z6�	nn��= �;r�#]���d���Oaub5x���s5����2�䬦���b�~xj�{m�^����-sKz�F�c�WnM�E[-���9y/6�X��+F˞�2FZ~�]��h�(�Ƕ��]�r}�žV�ab>ql�Vj;��6o	�V�"�`�`�z��jA	��u8���[�����A���^�~�tW��
_��l�R�V��ҁY�� �TE_��?���,fOc���?�(sf��z4\�C f�Up��8���Ym��/s[�� `�6;��[�u�2�,�&���d\bvf��%����M#ۭ�#kAߨ�O�\�	D�g�+Xs�ja��F��Uʢz�>CSm��1�m>ϋǡ���M�9�s%qb8o¡�ý-J�щP8]�9��"S[x��\e��G�#-�B15��̓P��HYk�_V;���V�|���(|�&�"����&�s��~��U"d������쨑s��������SC�`@�Q.>�|OY��͌�{�s��pk+�0����8i�׏�.6�)۹�ӻ�A�~���� YS�EǫY�#b����l���F�y�&�^O�i��Ỻ�v��]C�� y��(����5��4k�@����/הd�/F�!�}�/UA	\�>��;�a��B�KV02�/��ǥ�L��Z�87��U:����L���Q5�(%/�g,�t(�-���>��!�/Խ�a��l��\<D��N���}����xT��f�J��#�4/�;f�^��x�@/p~�	]9Y�>��B!b�N4Oo���	��t�خ��l���Ƕ�q��!j�/�:c��ZAə�0h��f��/�����9��<���U(Y��j��;���C����z���R��N�v����C.�STf4����޿��K�}�v�O�5�^8u����*O��|8�u��X��g��I6%���"��
��4���D�Q|��rl.����r�������5f|�ǌ�L���<4%[�,؟�ψntn� �[:f�̟�)��pN;��{����W����Lt�4��ќD����� S�z!�*tE�wb7+��5�Mvd6	g������`z�	%���g{6TK��^��e s'0�~���esfZ���y��j�\G2pVj�e����r�C�}�rwR�������=�����)���{c%��f"fT��wTP"Gh�8��xjΜk
dsm)�7v̓]�*zrA���}O�#KP��|@O�i��j�]�o`�+1��-J��y/#�4m^,��ҥmN8P�^�ia�w*ն��1�K���~���wS7&��8�oG(�����A�\���Y�-���-�/��x���t�AR��n_�ch�'p��x�C\b�Ͱ"����)F��wC�$�yZ6Er)��ְ��	&�.��]h�����W�9J�1TVL�żOFR��\��8�S5�A*�r�^t�J��{�C�"{����3�O����C`�Ό��3��A[���3�X�y�ܿ3�r+!V2��|�~�-ɐ���`߹�A���N�-�-�7�&���鎼n8��?��ޭ�����c[�R�d�^���W�5
�����3��W�	;ܙ��+ֲ����a]"������i	��g)jB��Vm� ��P��[��BR�I�R��=<�|�N#�������,����G,��-�}�IT(�B!(_���dl7�V�٤�<�w�V#���.��P$V^]e{�u�Ea%n QJZ侨�v�I�Sě.�m7!Ok�J�q�x:�k�S��iٗ+��ykWy��g�}�l�N���X�Җt�Ę�(7��Z�@'_F�.�_���5�^���j�w��?#�m�O.���.���=7V����s�4��NEw�~���s0v�����*7�SbPR~
g.�)�`ƴ8d9��[F�`!yR�a����7=7]ة#q�K��$d�o\i��O�#�u����ںwXb�w$(d��ؽ+��24:zLc����7U�mWX�3g�
���Mr��w�` ��$��3��۝��\~��pT��Q�j��M��-�j�
�}��i�2��~�|��لC �(��(Sz=%���ζ2�z��n6�
A����^����<Q��M�-ē0����0�\V�x��H�'��]I~Jt�]����_��R�&Ƽ)�k]v�EC蓍�������;w(��8�A�2����Ꞩ����?�,2rw�Q��m��R�E{�6�@š8��)[2��\`h>mޫ���L"l�࿨\�Wvl°��	�T���E�F�l�r�D��Y��&i���z��a���ˡ��z��B)>�q�c�y����#�.\ ��n���qp�����}:�5"�w J�R�(,Gt���p%%����C�U<b>�=R��u����~z�?�ޚ*G8"M����h���(�����"��TQR�tl�wT0���jn�z��W�
��Jc%�K�v�p'��O�m͗��\��ۆ�g>�G.�h��$c)A�ٍ��jJ9")S���h�#�-n>�,����~�V%.���P|�Uֻa!�9����!�Ó'�J���sF�jV3����I]�}K\u-U ɍ�^�����+~O�V�P\��BJ�O�r�d�:=�@���(�<F:{bh��<ԧ�O@�I�SR�Z�j�v��
U^\/"��<_�O�^�F��q��z %�J��&�:�W8�ϖ�����IW�L��F�qi[9�1#/�[� ���+����p�?���	�'w.�ȡD:��ՃoH�n� ���u,�07v�~ٟ��)�o�P�����u���
���x�P�+Q��.
��,�j��~ۧ鰒�N������Dǿ,�)�j-����Mw��^D[ؗ���/~�z^�?�n��rG��?����PE9j�ht�՚O��{� ~Gb�9�>c�1�V��sX��3�Ю+��h���by�[�������31���D>�vOo�Rǆ8�N�����m��������&/��#�������T�����w6,������j���jfp}�p*+��6sV�OT����3+�cL�������/�Z�BюH�
��x�i1�Z`[`���p�aP�\��*	��	h������3O!���dy>:;뚟�B�,zcv�q��T͚Ӡ�l��z7C)�c+M�%@�0j<��'���`����m�r2ؙhϴ��E����|������"D;K��V��`K��2$*���������_����˻ӂ�#9S}᡿*�+m���0�+��C7�|��sr�A3�R5O-\q"��J!��yJN7o�,�[�os ~����0oq�)��D*�j2��N�'����ȅm ���n'��"�
�!����N*�����<�j�+�[�vH=��9�$���D���y�r�k�Ȯ"Tp�]��aO�<�y�h�+��@�-MHqp
�#�`c�z,������J��������00Q�u�� �J�eV���v�����(Q?\�"�&���5決PA}.vμ�$� _�L�|��:�t��<�f����p-mn�C5,/���
��|�Autf�Ƽ`��%���V��e�?�t�(��s�c�A$��/G6��q�(�6]G��
��O����߃�dC�!&�������������I{�D79.&��@�(X�r�d�����h���O��(�<G�}昐��ێ��*ҋ���oN��[���r���+�,x��'�%C��qo��}dK�����xI|�P4Qp*����q�v�/�'p?�ʵ�#*�mO�R!�zw��,�^R��,@�KcD��K@yU�f�Q�[����`$_)C�����|�Rʹ�-Q�R�s���<�lHQT}e��uJ#@�Jy7&�sʪڝ8!�}:��_�����W|lv����ʗ��Y;�"t����]��g���χ��E���4��M��Q��Y�Z<��qn����p�l;���R	���8�,�{�N�V����AN����+O�W�S��&y��O8焆2�'�C����JPU���>$m.AL?nUScT��zx���!.�Sb(1=���U:mdĿ��h��q��D��rz�87�����k�l��Ղ7ָ߃x_݈1�(�cx����*�M�9!���-��_\�'<��#�枍)l�sG�)
-�[c�����Z�u��SֹĶ���C�ы,���l��V�t��F%�J�O]�0
';Dz��/K�)�
��r��ɖS<��}5� 0���*\�k*�b��!��Fn��5G�����v���͙�#6#'-m�J�ǅO;����E����p��J{�U���*���U��#�R�8����l�$7�&�o?�����L�[���#>!>�4�������� �"Ŷm��Brt/�M�t��D�[i�S��H��n辏�'*Ѻ���]c7,g%���e�nf��>�j�v	|�4��v�2�Gx�I,�bDyi�RP�9��ݣ��.���s1�=*��֘�.s����0M�&	�1>f	P���t��Hs�yW�>ǽ`kQ�Θ��.��h�KbƹeK6 g�����l{����<[b� ��V;"p�3��
,��k����QVbI#�е��i�6��6N��0����mN�:�jf�>�;C�N_��=��e�ȗ��z/Fs��W'�T���x�摗A��I��N�Î���z4�;�b">��@G�P��R:�����.�Rމ��^ѧU���RI"�k՜�{�ɗP��)�h3�Z��h1r'�"ݏ�ř�g���0dH|32�^�c��^�E%�1�=�qp�T��UW�j��isat�6�R:9�Mk��E��@��#[�*{#�쫿�?y��5���s�3Y���[�<�Qn徚@��+�1a�`��cb����Y/>3�U��m���2��]�+�%��KI��lϱ��x�t6U��.GB>�+r���_f������=�'�֜�.A�-��;��![�N}��t�x�%�Vq�S��`��SIQ}Cla��Ś]SQ1o�!�n��FK��S�W�p�˱t�T&���!���L��iNXa���Qw���+H�phbZ
U�F�X7���dR1l{q�Ŋ{5�ˊ���x5����Ci�� ]��h��M��Ff=�Jf댫t��d�ʹ��B�ϸQ�BL��;8';�s�T��#N�t��㉥/�B�'p�����˝J��E��������7S�x���k�u۞bFo�=���@�i7p؉0`Ӷ��n|�p���>i=�m"TJ:����H4}ǩ���-���6�ɂ�'`�2���*��4BD����<d	�ݴ�e���嬘 �D�����ZwF�F��������p��*J�Ռ��mA;F,O��~�#�8�Z�Y�s�b�r�G�?�)��\�'�V�9��L�I6&�� �@������\o;[��PD�;X"�:!}���}�-�/.z�ĝ-7o��oYrd�s����Y�h���gd�y���g�HnS���nH�F�Nҭ��Q��s
<.vЭ����FS�x���B���3c��Y�Ҷ7����b�z�g2�N4m����a*Z�p=�����H��_��ɫ3+�T)Vn�Q�tz����z;B	u���̥)L��V�r�@�ꈳ8s2�d���(C������� ����f^R'��8�xz�[��QQ�Zꄶٞ��_u�FŅ�-t;�^{�P?{�R��6����������<*�	M�=)M������\�h��d[��q�_h�#l����e`�����f%��ޙ�"A*<�!&�s�%�h�-S(��>x9>�
�n�,e�Cn�v�RǱ_���Us�r��>��O��n2=��[;>��uג3�����w��z�7Jg���s����(�*�m_,�'!K'&�ƨ���z��K��pX߾*`!�IIo.6���P���2'6v�1~�eYd�#@}���
�v{
v�PA,W�
�a"CT��vg���t`P���O�	|�"U���sd͵Ip`�V(���.	Ul9 jXe\����~����S0��Q�^�2��[S��S��+]��@��꾕d��#?:�|�ms��z���8�\Q^HgǛ�`V�}�s;�/�G5�+L�_�,�
����`�qp-]�������6&��Lq�_�x�Pjs�����tJo�o��^h�F�-5�X��ӭ  ��O��d{�ewA�����)lbs�#���P�:na��Հrd�A��c�̃�6�l�*X�W�-���|��z|�l(��tS�����p[@�������K�T�����6�>(t�^����J�q��BE�o� �=����MJ��Ȯr�B�-��������&�f�y:�._��y�(��I�أ�i�_�)�b�c���3!yp�>t��s�&#_���TX�nx"�=��+�}"�ϧ���ق�(]H��ZL�I��E*v���q���ϝ�M�a�?稟��"�i}�F�͘�*vd������[@�Mh��m��4��ަo~�e���a�a�H,���	e^.��g�<i᧡��3�8.�� 6S��
�� ���*t�n�����`>�L���=y���pײ�Ɩ�Q4ۈS��|��
���c��#sO(/'ңAjv}�bw�����7﮶{/>�yՠ,�7w�j���O 
�+��������g[A7��Y�� �n����G�Y1�#g���*n���d�O{1�A����z�<���x�JV�h]t�yko�ҕܝ��_�t�t^�3}��@[]&Pe�(��m@����_>ZD^�|���-��u'��$��H⓸-���7�{5b\�}	�V��v�0jF��O0[
}"��E@��r���|�cGs�n)�^���CT஘p����
��ac����6~3��E�=%x����'ՕN�ƕqt&��U��@���>FM�
Q(	�j������@�Z=|���+Y���p!�R~~`�֣yr��<O�K�e����x��%e�
��rѿz}޶���k�ɇ��/�od�z+H��X��R��x?{��w�L���$���z�pmz�58F���I��AY�����
�HKp% ���Q>c9_�g݄�3t�u:���U�|���|�ZXg�UQ�K�C8W�%���8�ǩ��]^:CNxxq·�ޟ>ᐇ��o�K���}1Gm�{����cn���ؐ��ݞ��zy��K1C��/;�F�̰J����H��+` ziA@�[�AKw�{��"C:���jg�x� �Y�r�v�^�W�@��(�Z�P𝸯���k�e*����3����'���OIV����1Te�O5������C��)�! �=\E�f��~�2�F{��1ũ^6 �x^��1�,S�n;���`�/o�Ͷ8k��<P_mmXFu�M�k|VAI"B��rf����d�J������l��@Z󆞲�"�wT���j����C���`�E �.���0��s��\֔�2�xZ0�3����[��>؇>t�X_l#A�Y�HF�ӝ/6��'��s(���zB�{���=�Q��%��oA��0Y�Z��E�� ˁe�:�Sq�� �����_W�h�9/�Xy�l:���p�JShC�W{���Sq�LgS�o<�N<7i�+�����;�azg(���G��r��q��k��pD���ͳ}w��sAf��9���ж58�فzFl�1��!���u������+�]Z���Փ��$yӰ�I)̵?&�Z�"YE%6<�0�v��ѠO���^������^��R�p����w�I���]3��x�H]�v�R]��^8*7�����4����-������A'D����C�(�G����$6�#�zXW��[�Y�j�D�.J��-�X���.qh�Tᅀ`=n�ޱ$���� �Vmy�0n0{�B~x-�
8�ħ0�7�	�E�¸h��&��h���E�$Ņ_��v� !����L���5�(L��n�0� T�:��b���֯I�EJ�<�ZFJ��%ݖXw�^��TV��QO`�I� <�>1W�AD83jA�4��֣ɷ9���^5G�j����K���Mވd�@T�"�� d5����N����p�S�y�+_yx�j���]=�Q�F�C�	�s��I�QX���r66�z� ��M�wr.��Jn3R��ElsC� e��g�d?����q3���M�<��MI�UkZМ+���t/�/�C����q�5��d��\ 9��L��� ���� ��k�^�@.�8"����c؄��l��V�A�fQ�����6���E��qBh�ϦuϜ���6����!�Þ^&�3z '��lt
q��&����m�LOq�!�I���SD|��n����imGS�~�+��N�WW#��v�Ppq~V�p��ɡ�kU��UPNYD��Q�� ��8P(���iec����u'�iI,Z��R�a���$�-�9�?���%�,Z���4����=�p��-Z8����@�x�I}�����;�n�dQ��{.g�ޛ��&��t*݅�DZ}QNh�U��[���K�34��]3��ei>R�^��N�{x���M;M��K���F�9�AL�ch�N�iA�B���N� ��~#���';i(~z��ɼa����c��"y畮�t�*���`K2˴�4��%�Z.�/'��C����!�[-<F��7���?0������w�`�ty1l�5�lk=���&x	�~qer�g7������y��ChYM���6���V�3F_�¥��X
�>����I��cA^rP��:�#�U��r������L����*��[���#�;u��UZ���4U��/0� K?�,O�J���+c���0����;֮AXk�����!O�Y�������ݭL� ��'\a�21O��{Vo�c&�sBp�"Ԏ�[O������O����hg3��)�?��2�l�N�V�9�}B�X|��6|`�i���X��g��>����M2����p�N�^n�a�G�@1l�@6�������%��JB	��;��X*��-O%���k��-4�;1G�k��7d� ��]Wn�sˏ��s��q{h,�����q) :ˣ�H�)h&xņ68�F�Ń��w튣��E�mf�e�uhc=q����D��,U4�܃;M6��C��N��g��K��xI�E��gn��V�Z(?̃"6�y�(c~����,}-E�#�X���'��'J���&.d�����hoz�z�}Hn��!��zPD�����N�;!���q}48`�^�c��?���Ct��z�)�ƃ���;9ҋ��"l���3ѵ�Bq�dq@RLC5�ף��
4�t��g���}���+wp-bp�x��)�^��I���9yi�J��aeUO���h��n��n\�m�P�[^��e�}~�m�H|���3��X�N!w
i}5T���6OP��'Z���jiۧ���O���ȡ�ڈSv������P;.���	�����;��p��W+&���QT���=;�����'9چP�ʮހ{/]�g��	��Y>��Ï�|=©��&���%�%�/5�� UN�n����~�[I;ש��C��,�V��e�y8�B�hq���9c��q�����b����w���-�X��E�jb߽�U}W����O�e��ZX
��뤗h��h�Wʶ3�����9 _Z��m: ��	ҁ��0�g8��u{���'�6M6��,���/m	�%ԱdY,�1z�hP�כ@�m�v�����������&yn2���t�=B+����Q���DF��Җ���C?c�p_>���ƝnL
�\�6��d��h�����ӫ��g�����h��]P]/oF�lQ*����/c�Ă��ؠ�E#�j�S0�kz:���b|Ï���Y�4���ϖ���K��&�٫�zM�TJ�s���}�&j�E��>%����Ama<I����0
��;�8��sY:5�oՂ���M�`(	/�5��L rvf�GW��(.�cnL~�l$��#>��B�^CeC�ÞP+�7L?x%�4�Z�YcY��{��B���=�x�40�
EB� ���F���
_Z��?פmi�p���~@���JJE�W�X�%����8"���*���S�>���Y��ʡ	|aC�pK$hDA�ǉ��S��\�D<=Q#�8�!e-Rb���y��œ�I�Gx}Xx��~�O o�hO�`êh�r��O��M߻x+������ �`l$	�p�|��F��I�S�lߞ"���`y��w� ���Wy�D�f�L���� 阗�c3{u�;(�^����^�G����$-K� mot�"Ѕ��$��=ۀ(����j��ra/�Z�����<5L���8�	:�v�HeR]C|����IA�S=.)�(Ss9�X�������ȩ=�C��R�\X����V
�U��w��m�k!�Uw��\Jx��zC���'uY?�Y1��)���8��ۊ ��S���l�/7]O���M�(���K�R�g��T��䬳�����l�d�S��H�q*ss�i��e�W��kiHc�yk#��FԼ#�1����5!(����r癎���6qM�~)h?{;�	�b���И��b2�KeE�ß:�ЦNi��@94���ZQ1/���b��B-��LTťB�.�2�q#�PtGN��,�eG�dU��Jev!D���h���C�����|�r����(��)
�e�K�|�Ԕ:�:w}N���*�&�iƛ���G�O����ȵ���t�\��uQ�إ�G���<_f��Y����!Λ[�4-$���9�N��m�'��뗻�z��Y���Bh,��1*��A�ͪK.�?�k� �w���KfJ�P�.� �}܍C^yu.ܷ�@�ھ�ZE�,��~��#X��u!]�����%a9;[`�Q���!0X��G{ �%��9�
�S/��4�ia�d�b�R%:��B�U�m��I�JSF�'��D�����|h7j ����7������~��ת3"Տb[5���f"�����`<	�UH��Ȗ����F���m�p�t�_	�Dtüs/��O��������;H>�=-ݜ6���` ��A��c���vyu�o-�������m�7����s���	���H̵!E\տ��D��{#�o_�����$T��UtDD����id�f�������&&Lz�tt6�����04eu,�E��"i{-�Qb���e@^�E��g�z=����\3�
"��P.�� <��A���ab*h,\H���_%��;n>Tx��M,tFs^N�������`-��4��7ǅf�m5�~�DtN�ژI��Z]L�������^Δgހ���������2��:c+k��(C�S�R)��=o��@��#��;R�PӉ�����h��q��!X*3	�Xi�I��'A���1wj�	ư��/� ђt��G��#�^*�)bo��ʠݼy>VY;��J���9�%y�pp �LѲ�n����oI}��Q��6�(u���J�ԙ���o踝S	8w@�f����0ͮ�c5�h����$۳D�JI��`~I���m��W����P�A��Iu�������\�k^�S���/�����{C�<�������d�k�������(�&��V�<��5Zėzr�b���r�[v��H�5݉�pZ�T%�z���~⤶u^�␖Ҕ~21֔>x��բ(_�b��9��z�!B̠�}rv���i�.A=�e�s8�A	i�����1%�i��6�k�(g�!�1� 5Df
�G=���#nu��ЧT0AL/p�&B*pwk��yqf�۝��r��t��s�S1�D%#s#�8쐶M���\���ԩ)LQbf/�2�IXOOt}��z�ÉZ��{�7�qQ�i�b��H�й��j�Ԟd�/���O����~s���4j/X$�kU�ұsO-�ܢ�vd�pr,_I�)�m޶�@-)�Ϧ�A�}�o� 3΄21�Q,��Ro]hP���a������C�oyܯѡ��-�q�q�h�y��%��(w�-<?}���
�X78r��ۚ��f ��p7�3]9�4r��C��30����Q�ɬ4��0�W",ʞ5)O5��YU��KM ��@L_��q�LȦ��&�/�7ځ"WP�6�k�C>�!��,�T�@��v}����ޘ���w��.�,��a��͈���Q�סP2�K�eh��$��O]�,�5vYW,^�&���JMw�sӎ���w{J�*	{���Gn*C�W�7 _Eh%Q����!��R������F#M�� ��{h<��h�!��ig���܁Q+��Rr��CI�K�	�;�x׳�'���ߣ��S�)Y�c��D�;��'��h�6��Z�'Q\��K{�I@�KJp��q<�0���%������N�r�fr�&��>!؝���H��a����9af��9��6��j] 5�%��դm��B&>eR�C!�N.F�����3��o/�@Y�# G��W���¶t��*��>M��%1�(�0֞?|��_.U����"����v �^��
 
�ӹ���JijY�N��:�*�:�E�4�%`W�qs�㯌��J���Π\:�U*���]����N׍)-3bnDZʖ0�uxv�P��!����C-8)����b>V�ShQ�`՞Xو	\�@��H�YBM.��w�P�T�啪(K��\���ޥ��������5/��e�i\�")��+zf��.l�ލ�8�(WB>)�>��b�9�?;���`mI�O�l2�Q�ˌ�z��v�0�L����A|l=��s�L'�u�3��t�L��TV��.���ZR��<�e;���<~��߶�r	���wV@ x��m@��J��M������U�m��zj�m�R�u>��{��f���~x�,�tY�g� �c��7�4��\��r������wYr��þ�|	�d�����c��x�����(�np�BYuy�m�-c一Z����Wߧ�3�sx$^0-�ɭB#��2��(�q��IW��Ac|�>�̻F�,��=x޳uQ!Ƿk��W�9T�䠞��7�y��6_!e�>���NTă�a��Z��x��4�S�>�3"B��?G�D�����u!�uS�²e��'@4����8^�Ãq�8�v�=��5zl�WLN��.� �А�����.��T�����{ץ�F�k��T�D�B�E\�)�&iWC"�0�Ӑ��)4�^��U�/'���!��i��:B�\bh��#��cB�hl�=���.^����U�R��iS1�Fsщ���&�g�ۮu���i��Tn�u�_}�j�)t��P=#�iK���_����w�k>�t�#��8�Z�L%��i͂h��t�`SEĹvL�Vxa�2*�;�-&s�y޺ﳫ��������H2H���f[N��`��^�� e_7 B�#�L���=Vq�1"�:��<II�j��V�P��=O��tք���_2�o��9:����Ґ�m�|�/�������|�U������
B[��l ��x����g{��������o�s���I��W+���6��5�Ԗ/8�pa��k�Ҧݼ<��.? A-	Lw�٘�y�����H��Q�k��(/�7L��4��&Ҵ*3�z:<i������)!�NIV*��\g�D :d���cN�kc����B�K�(!�F"�����>����+q�v:[P��[�Ou�V��eҡ
�]�0�ԝ�ͮ��2h��	����'h`R�Q�>�n��<��h2r�6�#���RP
����D��7�~��yW�dۓ��Q�Y�&L5#K�-k����)��
Ӑk������Th�.Ly��:[���e�'X����ؠ���"�#�r/���ϋ�ůnh��{D�뇄���y�sI+�{�����ȕ�Io�9��L(Os�k�t�n}��%�Y���͋
;��W/!Q��������$4�	����Mu�k"H�)#B��T��k���F+�[�P�ĳ�p��(��$@0�Z����/+�lp�1�YT����N>�O��16�^Ac�S�"�IX��Qg�2�>gx�� )�Rg���_x|��բ՝vf�l���S��g&j���Ļfhit�O���ޏ�d�hm�<Z�Z�?�c����v��Zk�t�<-�h宛_���l[8OZ��}�[R�ɰ �T�c�(&���� йy$��%�O��^ia�Y��f}��xf�������|[#�>�j�xT,�K��k ��z��M{_��¾j�JG�C�$�D�=�RB����Xޥ!�zӡ�?�:hq)ȎX$�B� �|�@9��78����޽���,��oH��?z��
�K2�r�ӭ�Ěf~�_�vK�{'�emY*����&��{���R��'��=+��
r���>�e��D8A�g���F�a�Z�Բ��mN�Kv�\-� �ݲ@d�E' �7t�x.փOB�<{M�Sj�v�sVO|V\⑃1��l�̢�*֫fl,�9��!'S<I�-����r��	=#�
PQ�����K̓�����]ޓ�f�_��?���vVy�o�ш	=钾���8�#	bzp�=��
��4z�~�5Ld�<3[![�[c�������|Th�N\��?�݀*��������N��}nMXS�%*��e�OQBW�i�%���qh��G˙E�$9i��r��*12E�G���'^��Icr�N��3� ^8L�=2�Wwi��9q- ��UQ��m�Ŀn��T�T�9�]y�W���qN��D���o�y�����Q�x>9�Y�)��3�Յ��y��2�*�hvb���A�I)�S
��>-���5!s�Fu��ק���I���?^[q���y��`���Mq�~�x�� Ew�b��&� ��L��6���i$�.t���L�B������>|@�H���1.��&��G�D��kѷk	��z�qUu0=Ά�H��\;��-q�a�I}�FS�M�W���8�tJ�����|��vC��Do�:ٌ?�CP���R��`I���ۤ!�4S�Ɲ���
@c�
Ou-�Xf�c��,�d3�A��������I�,�.A�ս'/tT�I���j]yW#��?;�,�]W!�U�ZE��&ٿ�5;$1�{�=�H���%�b}����I��������ہ������e-�AZr��:�Q�HN��2�CK���1(R�n�Gk����`V "#�l����J��C�aC�a:�.��oe��CHO1�K�q���aT�j:�pl��<.	=����l$�[�q��<�GT��U#j+f�4�ΘE���1͊�E!2L�@�7��`%�����wF��i���v.8L|��7���c(��<�)������ny���!�H�7�xq
k�U��E�8U�@M��|�ul8��� J2�8�!�T.�E?�