-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZbUy15G9PHkJw7+oQZtxHt4gFf0f1G2nA6vO6mX6VluSc8Fad3akhF8Cy3kyMCnba1CH5PIpvO1s
I+AjKKPCSsWUJQJ2muiiOJkLDtcdYNgm5DjOWBqWmvly0xIRWpoTnvG/sZo/i3mLFhFaEhcqFIJF
xVkSta9evCkU4Wu7hhVE2AabPYzoQbJ3MEIO66gJhmdeBJx6LWMoIDvpkuRZfLb9Ugm9ghXNiCLQ
Ed4mTudbqguSDDJ7zv9LqZ1zoJ5jMzJ6mUO550vUexNmwa7bUP5CL8Q0Tr9QpD2R/u4RT3FiTT75
uaGMYsXnLatTq900nlYXYQ99XB8jJ1WLkz/Blw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9760)
`protect data_block
FKhW9OKMWv1vCKEngszlZlNoY8d8uE4hR99g+uUCDBGBKkWbCOXJ4B2duC0T5zCDf7W+xND5vw92
/MKYE/kBr1TTrKzUCCshWr9e3WcZkSp9qhMeulCXY9rlPydX80fHq3fM5+3IaTfTxt2VzEwpyPUN
+3O127zNcIIlsA+klsDuwgZJdauQUM0uuk7Xk87j/bWLA8UYgMOQ9q3YV/SZtOB/QSdIR1gGQzuD
oEs6jlME8zpUDQRHt9smQdqsyhNLWIT+NoF9lshZr0FQEZDOkQMMdAK0w/mau9WO+qMM/kevQ3cu
ILqTS6d0BNSRuJzywyewcKQ1WNsdSk81rG5mNhsKJeL/R1dTILxFSIpTPLAD3I0hSksp18CLXIUA
UD1H09oQDKpwrP5fuKAFQP0+MKUt2cMxRl9iC1D6LQrcHczGIFk8aozx6Dbpfwtx2ThLBc6I0ZB3
RclzGhfO0lPnjJgFlT9csT6y0djHEYdL8P0f1ALevGsPUbqgjv2I70UWoAs3uf8xsfv1xQJAY68u
ikbvGG4EMliwx14kb6hht3Z3ObEucGaWmI2g9JlyNcbCAR7ks6mCPHdU3kVspjJ0LYuxOd+oTBZU
k16CS+UIaqDnsiT0e1465lrocYRpMGtwdaB05l+RFEg99ib5LMAfhV5nkLrMG/8VnRTOhRmgPor/
VLcnctgj3ytsdhQ7ML5zc0E7TtP+BH5ko7LKiXWlVhnAvEBWl6k6SAMvI4M0P9syG0/Gut4AXLc3
uiTXKtiZrhZ55Cvfz+6QReKWRb8E5aK6j1Yjr7vTBRpYe4rFbgmue8dNpuTWCxhswkQgy9I8UcHs
tsTBhWEkD2rs/xnJ01t1mk30gdxeljNaWWWd8WijVsdlssIgGYGJvFqEZJ6c44fwd+TUWh1xzCbr
T/yIGLQwkx054qQihFpUOsoBQwIl5SxIYv0oPLe4360sa2vr+YY1ezzVp9NzGp9lCl0zCjiEUqXt
KcknaVdGcmOLbNVMYDP0c4myUZJ51Dw+CJE/o4xuuUpabTbyvvIl/uq7sKrSqhZAUqduCWwSIIyo
vDcBr989Q08Fsnjeptc35G3JqL9bxlqGng1kx2I807uWZufJTikK2p/4g+F2bIRhOzKIGhO58Jcp
ZJkE6iyYMmjIUBjbIcweZ4E2LGdDYhWWSbYX0KXFacwrMm4yHBeeXRqYMiCNYaIE/Xhp6MDOL4cR
a5Q8j6NlWH7Jzt5WuVXX8+7S+W/d/FIoBs7vZjr3HFZ7FY1XMhKPXLovK0V3zfDmuGfnlvPReN7n
rhnKpEdBxl7UoLQI54TND2oHv/1sarHvlOPN3O4usuJRjuNIMaS/5v/GnCdpXW/qDdhk7uDnWpTg
KshbtSf32WC3dNxzimlu4QlwIG+F8pEWKWle9Mg/5vKQLoLuIeYhHzfZ1zCqF1JyJfZVl0OiGH87
iBMmeCtaZdKi62gyXcahq2nXjRA4FNrANh+c0AhWh3YChzyul5pMxpEjhBtETsPCzNsA4/IqJ/0m
mqqdz5j9X0qM9jIA7OSub4tfgy3i0gQoktC4mTsbmf7QyxXSExr/4HvkYF41CHpPflKihQVmHUu9
TVE2UEVxrzXSegoww87PaluvPCDlgxG5K9RmIMY/MJiV/YpC5PdwBH2EujSQ2cR+sfxxKiU/tmWk
NptoF1qiEaz3kHdHSkKRD3oF8yDmwIBd0RsxJCN4xGc0N1MZHp5XPqKE1j5QBRen2kjcH4sCYArc
Uqv4zzsIrxrDHZUjvZATy5lEY0oyUxEcJmguOqG8Xz1xOUSon+w9nB7YVF7pbtfp7uV33R8wMnXh
QM/3ytHYG/4TyCj1NptSkZ/KQsGyMbZUQAEhsgJn0BqpcSSEYpWW/dsQckqyHAYPPD5Kf4NoDffU
O7RCtzM5eGQXVfBzmZqC2/6LQTPTtXxJMK2jaG+ibJN/7SqRjRY3kcRjJw0k2KpOfarfsoLIyI1A
IZlPAwStpFPFUqFza/2KgHumlkq4xuj1Z8QNVuenRA4Qpu71trRHKnVZ8KCoTw/8PTpaZ7ElIt6U
Rs9+R7j0xacynzkLuijlJq3vWnIC66ypR/OAHCMNKCxKhAx3bS7EmzEYj7GTWFlr8Q4dqK6QLNFA
a/J5nHoi/YGRt8Gt5ZD0EZwrgMQG9FofWD4HYB+X2PzhJ0GSNIVT/qU+NccKIYN45uokLKFv0mVf
0OiTRXqQcKDALqIBRZFqUtJDqR5qYl6qv409MvOgeUWbDs8NFIajWkjZgagopxdgE2kM33N8DikS
NzPYY5FOeFBFHl/pkUIJAoS+Hp25q/jM8vsL5xQf7ep3wVhUPkOcRGm63ei45OKgxnC1M758sLmS
aNSKd/fHqRl8eAdV3VpicBGC4BowIx7qbDTpPeGjRetxjZO1K6LBASbc2s40ppJW+kg6bgZi89Q8
V4LQTH4egt57HuYb9CzE7YRY91YAADCMAgDws7J7lM5R6iFLBRvBoJfjwh2dH0OoKZPDUTHls961
SjnLhNV3urzhF4gGCWrAED0DHJbGGm+s37pug4d8TrFTumaYq6JnDbpSXgD7HAZNEwxK0HK6WJw+
/B6SDq6kJJS02jHNdcZ7SdLLYA8yu2SSA44gIZ2KT2rrsx4G5GfMdgKR5EML7zH2Zgm+S3XBj+vn
RpfxeEyPi0bPurv3Vm/5ubynOe6Dwfeb/nP45qvRyYAXLvWjiW7ucscj5wdq0P52nAnwiPiDHYiH
nNP9CEcFTmJWCK+WXB/NdDQoqrtG2pjTHHD2OasmoGVfIWLYgwGF3FYxGtzCZr8jZ7VUmFZhNQau
ZelPSnTX0dgosL9ID1B690JWY6RLdkKcZPzQ4RveVVb3PWbFoQqdI+hoFBuYUMqA6XWXsdXnPygn
zoYac0txRxPZINQwqI3cHr2QeQp+wv9h2h63WzvGLpiqxHGVHUaIyv0b+GlVTQWkiZf2xBdFwhKW
NuwBjldRXx5Jzfg7PUbFW+cDHRBe3SqOZwoUqcLzbeO6VuvxlHKlNGv7azNVbYRh6hWre0vwoQHC
4ESLtuXJ417vvtPkYF28KJcNqjSo3em7HmmPN+nYhZ8UiBjgMkxMuSm+BGhTpcCTslw4OoeeMqiv
Ru5eInIPNZiORF3uFyE9yTqzrqil9047zi9QhZhddWBmi9uuuyTFaOzstCkUzWhTyB6YVTji0u/i
TqIQrtErE+kMPSaDsbZRLjxesugeY7jMg46mLnF2kEK1lm4UV6pPHRvbn1Q5yAMpPZmGF89woCQt
GiMJ4bjICeQsgi16VMcNHfTLEWy7rLvD5pKr6ZM5S8JMghfdGa5RjBiwPx9CncH9cELo4kHhkg3J
dcrn7xuUH06B3mTcK34QW50qDkWTVbYe/B6QU7Ix2QyB+TuAZPkwxa7/P7FZcd3KIqR4+YkHDa90
4QZQvZM1jS68FVcsnx3jE4/hpVxItSdffFTBOgw6aIEQAWQ+SvyWBmydyWeTy6MpnQmIZmE88jEH
Ojzb73gr4qNxFnhdcX4zDLDS2q9aiMK3Xtk9ukTzvHDF6MwOMpsiyJEP1YMByUivqFs1LAbs7KkT
VTSO3k2mdtLxpM+cFWnXWBxPTzOHYrllEw0UaxDgAwX0hklOpNoRDibsJgfppNr2Kume4LSdPkI5
4KHqLLTPxUmQaZqfA2P79Bt9IljFpjEyE4fWmLPfzuzWikGIxAghAqJrfQMGwKvCjTKHZQxwv+y3
YwiTsMyRTCognOzpiDW/TMl5Rgqg+fLNfGsa3aGpx9e92DorzHfEIGt1122lH6w8FuCt44kqE9pV
uUGfgy5tL1q36X1yQp8chqsTnu2e/7gnY576YTaANgiamuG1d0tRxTxeSQZfA/cxU4jJ7I0Yg8OB
wnjvMhupKJUyKEtxc48qOGcWTqYXNNfF5VkTvVgjLPl6vYi9SuoKYc78+b6arqqzztG6KnlOE/pc
zSIs/K10kNJ+SZ+PWi1uquvY2lIRufxALtQBUDdnQXpXL93VtONQve/ZPQxIZkIPFVo4U1DFgWQ6
UmQ5Cl295dpWMfoIlZeQJRqRiJ0dzePDbZyrNatiR7i56KuD5qSz9LbfBrKFC4In8iAVv3yqZ/ON
u6gK0Oc/jYGx4LRU6zWod517rplEHj1+aJznw+7liAFa8KjphJ+FbSYlO/iGOK12QokY9Mqz7bdH
RRjiTYMPwLUk3QWUsfbyoALhOV5IImuWHGoiz96qKBW+bdnX5zBluOs0A4F6q65Vo+V9yG91HDjq
P/UK540wWFWt7/J9uPk5IXAfX9OMxq7qyUIV5danS+i1lPDem8zuE2imGugRI7dNjGRGlCP7dvrW
UnUDtNedfXJEESVq5uWLW4U0vOvtppHDz7UzAhHdK/sa5JlylHF3hTKM0zT2cLVwfQ4W+aeiUBfw
UNc/HGqAGOoqR0n9lar4uoa0m170Z9DcJ93jcPk9acjEy6k9YD81Hg6kd03FEGoGYB6axVNmw1GM
eJ8PBIC0XL2jeMj6spxQXlK/ucEkr95BuVwjz/1DZs9944Uj4AcdkekPyDzI/sCt9GYAL02mDEHi
e8me7h3lkYouaJH9wpnpR01SJdMN0Zylx5xFN8SQFLmqMIYDof2ovrW+s1I5nYyUwzKP+jSu6Ifh
sbaDLAXhPeZQjwxEe2FoD5Wu4SMmioRxV0GU4EMVfS2JjCpsin0K91BYIjugV5mBlyP7vlw3SGge
di3YCZeja+0KXp+hZOf1SgCo81lZjAHSX8DCxD6pPOJMmP5vf75/z6S5dgjy+I7y+m1qi26EsZtk
PujnV1WSj7/cfATV/DTGGfOEPXgvjbR8J8TUdbhtK5VihfZ//GUn4jS8U76ar5AF5BnIGeYPbXbZ
agu151GwNsgBTHIlINTOkBaDlFczrxXZutdmA0pvSognKBhkr3F7Tu36TjUi/1K+HCPapupTLOqH
KFTzIB6iJD63ZCZKRi27MSAbkRAIU+zg3wJDFFJLmzIyKGVWKtjbY3x3OxqzR/Z1QmfOwAufHghw
SiW9Jfwah/PMG5iuEbQLl0EP4jftqjtjI/TUQecsZwyPNwgkltJmxK8uC1egLYICtyj4lpWtBqVK
6G/sG7tmO2xeDbWt0HDeuwcrkd1R8jSXiBhM8tmXJ5EMdyiqwCqy9k5ff1vcVBnL/fCd921JGal/
uMNVVgXgJ82zfFx+Hq5T+58QJij7i0ZA5fejoJjJ4p4FA/MhiXt9w87XmvM35WEAc/LHfZ/a4PrC
adV8j8Dqadsr8wpPmYs0AauRfAHZq3DL6YrldEfoErR87Ama6S8vFtWlIzlgiq4HfgpLuceRKDPN
V5eHMf2IHIh0LNhIw8atLMGx44dmQ/X0ij5lybbEVmT/+F4ARdbJ+glwCUged6DKlp3dAHjMM3m5
z49Y5smil56rDdb9hhMV4jVTYSDJuUJxV4WXOf3gR5w8+JeDRpFKq+7o3bM8HAp3VoFlIz/FjgyS
wEYreiTvJ0iJ5T+pp1BL24bHzBLb+pHqwMSc3Hpzi4+TzRncEt4MicIdGvCeK528j+sCrrY/8XRF
cbLIAESUvReN3xtQV1Fh0ALjr3In4aUW2Qa/EwCn7h2KGPR+qvcl3Z2KSj4caXFqaG0kXYeE2FBy
iVi21urPyVUNwMYNskXIEjcB86c79eekOJO0V9pppZrQ4S0qU/QJMHfnIJ32uvXBeCwEAFM7PkOM
2lWZe0cOpzUjHkDo7TBiWBoyJYo60+KhFZpiWZn+fS6rHaGbrhSGAN55vjzEIjdXDBr1WU0VKEfD
qKd0Av2U5eqHD93FjL6SQoUb4iOxWwukfYLKKr3IzFcssvbke4MQLmfIey3dpH+RE5cJ5arsi1o/
exxF7pjqKBa8ojf/cAZcXPjsJdRoi0xcRMxim9CIkG85jahSNP5K8w+smDCC3hd0hyyTdNhz9AtE
jSoFntXMnmEwMnT3cWKmDb7bYw7Qnp/NpZAJPBZ79n6Zuhggr0D6cQ8/uSIwuNGvl40dWZ5amaOj
HuvXObFzXDVE5S9W46ccSQgygMRjndFBaxCfUAv4OOO33zPid5EaRWKYnOD2diw0S9UhA7pjxoTX
SI19cplQM65y+h6zkFnFlin+b+h3sSk+hDTkMgzW9BLyKp8q9QkB5AGMM/4dNUPPX6XcdfZ0qtWk
++6fE0s4bBha/FM4vm0cY3CTitcnfiNAMXdES6fDZ7is+bATpUWGjN6NmixjksTJ0VOLxwFGiw00
uWFj40DVMZsA2c/mtNza1E79RyalijY8erwObkCuXmiXBYFRecI5+puZ9h3xvnjFRXUi6EtpkKP+
TKTskpmTAzJ9WErxQduMONOG1xHu7070jp84h1O/g2+ZzAyLakMmNOkGXhaiIDd1PS5yd+hU6fTQ
2pqyjs828uQvfdPFa6GTTbiYLA8dPBHYW2nz5zrUnI/TTWHzHvwwRzbYSZmLz8fpG7DtVZkATIAr
B2aq/LGZn6hFdziEYFIufJjLh5+KrO3kR1QPKq80iX4h5+I0q/fi5B+gduRl5lIe6gX+XCq+rZL8
2Bcs7l9gr48zWsTttTSUvFpAB5BOAiAOpt29QfnJK34uS2ixcNwNCHRkoGmvPYC5oNs5E8TTzo8v
LHmEjCAPdo2ORZK+5Qw1TYZcS92DfQq7Ja07TzAjC7luAJT8TrOQy89S45RrAaLdtFPl9EaHZx9/
3ZReEubgFElmWAZe0yBXx+e7jUnUMOC/rZOanwKZW/aDXDU4/AOyFn0GuGi5XLmgQ7Wqhk9Jc46Q
//fvk1w9A4m6YV41qwf5Y66A5SKxcl6zDprF10gtHIh6P8Vg42J5nh2VxovV4DV0n/lWiG6VZ2rQ
8fCp3TlxqbFjhoq3S+sXz862huEiv70V/FQz7eMMOE305Iqj8qzE3Gkavd253KnOo6WDfQrYBvvI
VG7idg20a55qc+q/1C2hO6lfEYCM2Xw53dSiUI8COqd0OIRY4bxwlpP/oh0U3FNhIec3tJwprM0b
Q6+LBhB2rlgvE/cH41fpXpZIAUhLbRHvMQ0wzoSPquy+1Qbk511J6I/gZsto4hUfYDGntxVMuDbd
lBKgJqGeKxGdjEgQ4hMOlU0AQZfqpBeK70rC5775iEMZAVL8ArX+agr7VscyjH2V1ujYiOtv91Ix
C5a6heRJ8l0wVICqfWgm/HX+LjwOiZsemcsrQdIcOtO0XrXUEYhoumxaGuKh6IoDvX3BNQebDDTQ
i/zp1KnQcX0dhnT1dEl4uV/x9tXQnf95UpbEfXvJHffHio1ETdb7WvIdgZBGfntfZ2wFYy7jxG5l
F1zIY0oaaW81wXYX21hYGedI4+ZFt7N9G7mLcnuga6xh1gCMPBaXoiupBSnn2ix7wATM8Jg/JYSr
n6dOlUi3oHci8ApqaTpU+WZ0m/TuFjKl8xO5RFmfiB0A1QCE8tUyhz+qf0XQkioSueTPtuwkE/CF
pk+VGiyzD64i+/dRAuaqGibgk4peOMGP5pSNttCv2IZ8BeCzvn/FLCBOHe8FnRculRU7wT5hMqu7
bclV4owbJOCrx9S4nQ1XwskEYNu7UrhSDBdv+OsYZWl9tRpoohAUJ6+vN2xwLZ337g82vp1NSUsm
pE36/nHbSembYeTNHnidiPkVxuINlkN5MAB+VD+sM3qk4qu8W6qth0AsW3+oTmAR5u0/wM1194ez
pv8+WEoY8rTxv72lyhMilTaCZDnj9aNhJ6K2N660JKTYDf/DDvuDPDG0B8IJCEXvXwxlijcnA3iP
94NEG/FkyMuMVyglLGuyQU1Uw8OGiKpZ/mBl2n/ZH98gNul2OpVuczitYVmgFrtQR74VbHzGB8UI
bngkuyL6o783tmb67eaylhFrn7vqTU2ANcrOYFn6TnuhTScsz2u7cRagTQJbMPUzbc3ugfApHLLP
Z7i7qL7LLXP9+n9JIEMwHPn7djplTcDnHr1nbQE4jYbK6QCEEiQrV/kRyCS5A1ssscjRZMqyMiln
eUe5l+7kaTN964I+UebWR9i54jjfOpDz7CVH4Xt8qBuLUWbIe/vHblP+oyzq7+go/8Zla0qxnAKu
fwEF8xbIptOBT8PwTL2pg8SzF78DylVZlFlmUS7XueZHNPCJnE+8tLtZtNGn9AIc6fThrQZoqBMZ
fZqJ8UsHgKr1zwLg8CzLHLpLSy6XmbU2oAg3obnOxoyHbKiT2Wzt0iQJk2cmnUWjWGMXkKptsCiV
aa56Fi/Vtmn9RREg5h8JUzsopgKJnbxSFbLV5i+KMu8I7lOPutqzcgujy84UC82MWtWnkUgigLff
1ULljUkORGPxJjc6e2MjENK69xzRimm5JAcL8pDnqZ0VVJirhNHN63SUVRVporW7zd95AHHKfBxQ
SNO3orlQvCGCh3aRdWTaXgf7pTigIBdYFFf6AlsRc3yj46IXgv8EjgkRC0+fGNmWSsocpwi6Lu+R
dPGx9CNBD0/ZbY8C6gzoFJV14G+ZBLKjxott+Zf/ukxVclnOL3K+42dka+GHphtI6Y8QOsKsUUbM
+bHayFg1P8ImpEZmAE8BXDHHz+ru/oE5XPoXM6qXHcXO1Euld6N+5AnACUiN34y4Pv02bn4XCMmq
JLD2Gl//ObpB9YE8I+tTyjAT7vwQOCehI6vGl3ZIV9XFGxgnZZwE+cdFL3sMFbknQCDJ+/Vatf44
96LKuVHqyVKMrBjRuDrtCEP6fBIuT8gYVPoIcWpLlPHyhZNFzLMmP1opBJbb1egtfK7XtdEb2jXn
M+nfHsrPKTlpApldKelw2MONYKm7tA3V/Pa3Z6WzO9rwf3xMMAvEwqgMbdGAZSDCZsyxPmzq+K9Y
TYsM0cLtYSFow5lI7xK4wRkqxIl4ChHvENqk+ofit9neI9fDWTjeR/yi5IsprJEeeK/go8HlUr1e
iU5ErI32CpACZGGP8zNeaNaspiPN7m4nnqPGIn16EOxvI+Nr5KodtuV5WU+9AJXd+Obmt6phd06k
yU6b+eLiu5YM60bY0r+7V41eTh+gxnnDE8O6zXqb8SAMYVUlme3MRExSy+J5gcKgkoDoDhhAzjZf
uBHErthp0KqU5ivQ8ofb5S72Nu8LsR0xQoW0LQx/3hdBf0XtDGesPMfbHJceoJW1OuVUjbCJ6VCJ
+qZthUhhIWC4s64Vdi4ReFUUNIj4eQ0jTZsXLmPK8rhxe1k03KaLADhNwr1O1uJNEwCUk4KTRqtC
23d08NSZPXnxVFNr+snUoIhXrTykzAdzBoCn7Vt6IL2RdsOTP+ovbEn+Nhv1yG3je66+MRsP/HAp
RAdqsfAaAgxMsRV4YwIEccFxsOGnEYCZhcUVaEtQVnupJPDEwqDMaDYJ7MXs2yqxQihy3PuyA4zc
WHT9kCzw8x8Xb19YULxWZW0HRVBoydcd5nJZuRkgQWBR7TTDX2UE/mzLy4YMwQ9HEu58H9EF/aEu
4gPwV4Zh4+C6vCgL2Jsh9YuxMbcBhp9m1WwPxstir3VByrutQ2vgiOztLdmPTi1Akx6Je+vdPUzp
Gpt5iyWobFj827l/AykMOD0RllnpcuuIywDAg7dVfPxUxkLyTFT6ni5Yi9ATYKs+ZgPV4ZdKo0Z0
iUhbpkbELq8f8hTMfPhjjx13Z6+XbH4BJUHjEEEPzFRqwwH+3Wr9gNWnfhdLfnm9HrcKqVr59yr2
RO0n0mSMddvuasWFu/VuT1wgchy1hvlPh1mX4cLEDtDPg8vqjCQE0f8lp2DMABJqZj+m13Xw1xAQ
PXkYkvDFowQX+DwjhzQUMCDC1IsBAR/f7Wt5f+M3UxnqG1ZUOO9RdeTHy/6YGKsj7gKXIoKx4Y8X
a2yJYfkFUbw8SLnniybS2et1HdQHx2VvjgtNBr5TFVxg5CnHIkn4OY94PZ5TbECdbOvvSW4fqwqP
7aAPFXFx+7TEt4YF7D3/fYQEvVQnnQRTECI3kzk+sIux7JFcUQnbsfySCjnzL9DlAXf8Xp0oqfFK
cy+mZHm27B+6v19kgR6EDIwPm83DoQqlDpJqZa81TNiHUk50ahix2t3XC4uI1eBn2WyPws7rCmQS
VsWO31FYoQUi+6/pfCUVi1j0gZ7ejFosl1rvWkEfRvxocGM6d98mQg7Jpj9T5E6IS3Tn7Z0VfHZn
0HHzX2XaeJx7sNZF8+10C3AvAodGSQ8Y5W6pWJXMLOCfEqrVncA3D8/WhFviRzXzvpv9jVlCM9lN
08TFcdgp33dgFFgPWyqZ9aURwP0zLoHCHQ9zeAfRX12soZt+kuCxpgsf11F4BMihnBJBkcAD/Gzr
IUKbm6IfHF7I2u1jN7oUcwGZc0YUYvnx6tHuSTNb39i8IjEl4jxfJxZwRleR2FdCqjQpsaCfG6Vu
RX+UQ22UKyArS/SDxULnNyg8Re0qKuGOZeA2Fm/eNWNdaLBNiNcKIhnE0+r6XTRnRHrzdyDpEd3U
yaYlgQSRWY4RtvEKNz5tED6CslAlMDUWX0BxRFpb0Z5m/IT3ATWSyTHd66U0h2l4o/NdTuhNHYmS
lrbKkyim0stYuu3Lj6EHosuoiDklx9n3QrzwstqePJrScWUFivsoxNzxNmPe1r5CxtDiHUJt1ohv
FM2s8TYndKVWEwIVxC78PuIhcAEV8GyDNSsBh5a3Q7ct6V6iJs+hN6h9PpOUn4JxyK/KuESoWuXj
fE6dPy8b6LegqOKnBo1eIhgNjoROG/Wa9tV3/32d8yWQ/ev5gKhwNza7+D8xLbaQ2s2UCcaZ2Piq
1w093ORPDT8eE7vQsUJM3ItGjFoKZQgjB6do0CyKIPEtoezoKvXxlviBrvyqFSz026sCzdo154qP
JFoiQ7oKldds8M/PoImMD6illuuXfjwfwJTwKkH/qUL+y/k96pwF07KC7OGkHhPJ+XXS/kNQ6YRw
2UN3YlTmRnVT76Nfb2EizvtOVUuY8jp1FexaKjABXxYFRI/D05tBz8UihEeOgvi9PPq6fe+57CVR
9OHVIObEwhirFSbmlbWHEe+XvJwZLMQi3AmcclTX/uL9A6DRpVOeTuenUhzCniqUYdzFxSLavfPm
42ZdJj2s/EGBTm/06cvhChlVTV3RblxcOE0sjF1qdrqdK/VaGzXsIPT2At/5X+gIuJCqIG3bA3i4
w9pvaipxYMOIPI7vJCWIz1k+lTQk9crwxsRQczSeVQtjc+sbuyFwHWTtc7pFRXEzIyl0jGfkYque
8HLL4MdDpO8PCR7FiO+WIyaewWO8h7ZLNb2leg5nagUujbiNiPw+oVb86YFF4LT4xNAn6StQ1Wc/
IN2RiXdA5bEMni39vJYsipRuGmzRFHFkOES5WTou9UkZ5nOxApEPhtS0sTu8w/6SixYBK1UqmQWW
k0fvSNfl86Q02iRrajminqQDL/bSBAYBWB0o6HDS6aww90zgEwlp7x8SC31XV2lNEAqDbWd4GH8S
veUkqeFlQPWLRa4to88uhOhyIne+5ZTh7gCr7GWBuapbFKHgm1IhvpGsSalOB9Z9SUPVG/h8KSm/
vGMKlc8RrHHEGXvE+HuGBaK+naGc5KKaQKwk1fdjOE80xF8WAqCvMEXKzy7g17rAVJs3rivYxPI+
yS88p7HBBolPWSX+6uec5PN8CWfPYDlIMlN+J4Ys0amf/snX4v/ox9Rn9JjIJr7fgEyF1KVax1Ey
N1DIHgeaX6L/oxVB8pqYd3r5CZE6QpY2Cw+DlQqPYHxOtwgsTSisIToOVgIf6q+4/njo9LcZ8XYK
clf9VXxVoe3yhbG5Y9iasJodhIMFpqXmp2LJJ0Qeb6bZbgWsiWkxMwpEaKb8FJ3r0O5LgAoeMhso
wpio6z9cIIp3ZnHdEC7n9KmkKs2SZW59E/hqY2NBvnDWOExNcsudMHZlYWmZeTM6aIi0cjxD0fHn
t7Z6yiSZb7SVfd8R6TLpP7Dn526SnnPaexsR9YyTAhdNOahhPcSHjj+M9ecDAUbfacB6WztjygBN
n+EtBm7P7uytJsSjbqrq9HKDbpU5o0uFHpTY/4XAsnVJfg6NUkVweDvlxFtuX74ks01RN6mxpAK5
8f64fDzU4+9TahmP7s8NaedjRgx2Srw8Y6kHwAWv2PktULiaujTwSbQOD9Ssd0Jfu5D7QlA8fF/I
SSxdV+igF0mgMysHWEW7dOVpOQmfUZJSesNesjC1ZCNqqtzyG+0ma2Lcm4ayKg/pOm3ADme44fcV
EBiBOsy+bKuGNnIOt9+9EMcHUaDyUcG+qxE8O0ARNHBut/wiVhFUGiOfF5sQ14A358ZwQKttDmVb
4Q0ZfcEa6wK8CjsKP1NbANebLYN/TOfDxJbdpdCTjSs9Rb5Om0HAW7D5QYzxmUQ5dgoXMOmTqh5y
F0zHyvG1b+b+g4UguFLbFUz3e81Ue9nlxkc9lLlpTJxUH3wi1fOLe0Z8gEfW5gJpGyzNvKrzc+xo
BBhXeJnOutyfvOU7VgJwVKmE9c/BVtg6G0/X60f+C1FSzCUA65In11N92kmfFyXXY+QWedc13gwA
CMVyzEZEAkAjERLZacFk3spzFjpjFfoEmYDwRiyYtjugeN/K/KIwz5y6g8NFoRlVQkVZpd1eXVSq
RtJnbbHmGLura+d5n44nb+F16lG7cAQf3kudwGQmqwcJDbk9+qH9+g6Dmqhj/o9EHpppFBV/iFor
U8CHcQ8/Ym4lP9vTkNvjmDTlM1/RYM095WJc2WdUdqMQStKLhfW016qFIDegaqiKBeK3wFL1fAuI
q8C3lVviS3lCL52k2RbVYNXJWdUMMtW6ngpKaj2l01a+7m3Zpless0uOKgvbNqRXtf3FDzR8oKrh
FzlPVqSUQ3hwowZSdZNczPnEEoYh5K4DwU3wA8knHf2qGY6UnKFqm6erv1psbFV42AaA6Fz2Wi6p
HoqgfI82O6FoUaffSgN2RzGBCjVtic/NClFt8HPMXBhvAK6oIrUyFPz9btVKT3+oi3SJyknJhi6f
4MlcJnud8HIcP6kr9obWMKDQX8FQpDkHxMfL/smAu0/08NTO0C7NIjbOxup9LzOWwHgaF+atRFM0
6BqFCrVizIrULfKW8w==
`protect end_protected
