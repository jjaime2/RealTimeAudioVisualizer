-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
egM6z2pPmNX8fwmOJhxeTz2BppSLF0lcXuDqRenwNidyco+fPY5Cseq307Prm/noa8di05P7MEWH
h81/D9Au/Wnp6Jcu3POQ5aFcHWnObIyusMPXibY4MuseYkuTo0xC3h2iZOKsy4ha63IpGJzsWvt9
c8nIx1rlg66lx/OjRhI7Ce5AoaGhn2ROkl9r+OUTj1FEopE8VgtvkwzUgGUwo5gR18/lvncG+74t
OtRZ4nQt7PxmxZ2yAvPgOFmTODalvgz+BtiYh2WRWhVzhPXLVphg3/X0QkxXEjp81hj0hKKxleHT
riEzRS1kNeyLgB1qc+Gsl0uSYEH+nzsOTvP1bQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4656)
`protect data_block
ollc+8c+xLnr6WuMqp/4yYbdzo2j2KlaPp91Xm64eESTomn51Bfm77FBwXwGEKoDSvGYDLUZ3aSQ
ei2CmHVcjbzAJEZVQzJtJ+IP3JmnWeTqwrUa8T7yM7oAzFbRoYYEkzYS7tlwvGpCllQjOpAg2X+7
Lm3FOZivT/MXw7RLaWw6W7vbgbi3uiAV6JmUb+h/++SKAvGgR0FfoFrMEygNDwe59zSQGUeFjtuW
VoRK5NMjd+7V8aaHtsA+tC8qS5B/8FlbWAGknJYIejMaA03RBA7nAZ8pkHfY2xSb1AN8BB4raV7C
kaMLmWJ3nw/t3vCDsixy73y0H0eZeSgcR45fPJHN86ICdooaYfIHU814d57PikMEjUIh16LJ7+9i
7Uaw9p9cP0czDn6JCA9J+csuC1dD1WeBGr1kgJIEPuXhV1XLgu+2pK1JvW2fbTsSWvSZY7lv+rpg
DKSvk1yCz9B1hUBq6Gf7OJdt0PiiDg2+tIqZCn3YeNANRKJeterWuD9KjmJdIcJn/RJy35046nZQ
mH5QRf8/UxtXWTucAL4tcKbCcIKXJ7FjdI5YaNhj1MlyI9TV/UKOHzi5+3SM02hqIMqmdF94V0sT
YGXblmyigoQeho4mAU32b5N+Un9OXVfqa1DrTBh9v0xVz0wvMe67/x/u3cbPNSbYL9wEt42YCG6e
LmStXJ1sVr4N+0prAwQ46sbOH6ZtI07CN+rFJHlTEf5m48UXjeA5RguMeBd9OanYajOmpcd8ZlWS
crHjPBuKgZEblc1SQXxfkxuW0kAZc7ma+38tt7U7pB2wQSZKiXR7+TC1iuv8sQkH1nWhTwxrjV4U
Jt7kymLtYK4YA2GlflreKILtjVweZi+tkk+AFZGN/3jTBfl01APrIMP5XR+rKG6yvY99H/baTeTo
Nmq47oiPx6DJ8YWcSc6ePSt6n8E9TslNg+oVG1OWXmpwhcMKLSCfxHhCoLUGn7Lhxf5jggiu7nWS
S1ge17ZdD7XeDaMse5bSMWd+7oClXyrRYAC9xjD7XBzlfevs2GNAx2NKB2oFxqfu8vcT2sqq1QLr
dLvC+xlpdjTKTcgM4z1hBEo0mgobdmj5KzuddVdwMXH1M6yE8oxKBJ1yHx4G1+3SgToOc7IawGWW
mxTMCYCGDX6FNAvREkCrW3YcCkPMURzHsIlLwekKcwb8gaME2WAkjxrbc+458hkwalfkHWQkB4xa
he7jefyvtssXhxWsvT+8M255h6O+IgOMhZpYa0YRko2Psd0/y3M5gxJ2fWYHk8y+2PCJOwxW+VjA
F/ehiqBPYngqiGZQSWSRtidExWxyJ0NAqh2+MB5UaAgLj+plhR00+SNc9He0Jj/nMuIOq9cLy3RE
s1vSG5u/pLSpIYOhmsvsxEKGt9puL3rIfMFve703Z2l5GdRbbDDM+VgHhoNV9Qz0YeKmUifCLNGm
XdSe/9gmaJjEfxui0EKNpfm4u9t96V6dS8vVoSVhOovbGtowA+rIxqCK99oB4kfswSCySwITjjhz
pYEV76lkaquJdg8Kr2pUJQn7rL5rbLZbPJZ8DggE39RPoeVA19X0DgxEJPxlj06DIlimaj1ze1sF
IdZc848tHxDt7lrwWb+qKkHHYqv1RfNF+8SsWxHwCn3/CMaauH9GatKjtfjpleCLNNfcrQEyzUZ8
7eJLfg2p4dCdsbdHgVq5OX6hg2XdzaOeJlGQEKqS02biUiUQYnI11cynDJikhfoDgEylwA22SCrQ
9Me35H4FIvkh6KJZrsBPrcF02G9ay2W9MdHn2aue/g++3h1EMG2VAnt0fAZ52DGrSv9n/iDpOFLa
26nEJomxblwX/hsWD4sFOFkq7PJ3jTr4XGfy9nQUJHQbRL4SkOhrtV1m8r3f3LnieN0Qvbv8204j
zXmVMiKfHiW19LlmzlmFnPsGX29Ij9wH0Kt4pEYP2UJViL4EOwcB+8CDT7mx8ME76brP08jQUHXE
3RHFycmQf2dHZOUk+0G70okuLh3sYRtY6yjEO7kz/lOigiVLP8ThgfHqui3OWrIPz004qGy6iWRh
sTEeUb1l2XEvUCe5ieCPLAHLXaEATexkJypbhIxgprCOSpVRcprMOMEq1XpPQvzu/i6aK6jRwvSq
QM9Z1KEO2xALbECWs42TF08ieJ31SHYr0b91KIL/8FZ/CZS1cVyx2QQ7XJQPB2QCmSjj7RGnPLOm
DPvRhFYF+MPNc7M5pJwJOT/+qs0qyY+tK1eumh3Y4cOanEWKdItPj51PKCA8OB/oamfbNwrh2mXa
+ssgP1TSoUXvO7Cm/n+NkVi4VvKP2pYAOCGehkxEnfaoj7upM+cT/mo9JE6WvbrTzfPJzukRXcI0
hdRZNZxzU3U/H3esTp+ETysFWTTG6zNqNveB3BYCsvqeihk5Bo3Us1AYpshcV7JRYVMc2CvLYeLb
vk3kclFzvaeu7VBgEQW/xp2qY1r4CuN/KTDGlXK+UBYOiklHLEY+w3ld6gzga4PJVvRFW8uGlp6r
yOmLQnREGh2nGyO19ns+JYtUx4flkd3LkY0MMykpp3fw8szXbtrkg3RV7lGaZycXWEtWYLimK//0
nXLTETTam0GykUHtrWZTMn3EztQWqVkDS5hZ+2Nze2qPYpKYILKRcM4H90gpQe+XKP2H6AjJ8InP
EmzLdeUSrv8bSURw8zJLuLzVhCJFMCLwKPTn/DR+EMkV1ghpX7w7V/XGchtPoibTLweYvRVrjIf5
pR76bJLm/XbK5FRMGwq0EvwnMgn6eU9RH8Z9I+1BdtqbCTYrfADI9VTs6I+4rDTrlDofs8UIU9Tg
pgVRpV/oAs+3cy0FaP2lHW4+p8T3K7pQVgKnqrM+Kw9m2Zijtlm0wdCqbbIRWqMZz4odBW52js5M
lZBsVgtjpTLY+9gD9qLVCwagOwNtUI3Ut6OVKSQv9SqqBxbQP6U9Fypy57m2y3EJ5ZxNyGkAXIw1
L75bzko/pkxZD+WDOmzV0Fw1B6nXlE5/VE+VVLG0ST86RYeMuWpzmz1/xhWY9auVnbDSY6TE/szO
hLCG6W77TM8jSzqHqrWr5JiedQm65lycxEbC9caD1ulUnj0Ato0zmkmzCSGPaGxZbRNWI8LONUOZ
fwO9L8NNTM7hWelxROPDR2XQUzjtwpQJI0/XJzXswY+Wcz9Qz4uw7Z9RwlRflu9GyzcdS31He/iL
pJsBUdAPgngYOHeHJkDQZFrqtujdr7nwuzeMFiKHorijj1rCZseuL3ZQNYeNooo51lFeTFWPwKbH
bDNYpz5t3cAh7cycU64rA5j7w00uYo9+S5BJzw5h4ukqggu9Efvo7e4Z9BMgd7sGB/74oACVOuPz
je4ON259RofJlh624IveymosiBiFa0bNzZNjZSqXjKqPH5/Fq05mP/4R0QM5OspaFk0LZtofjjKY
lr78tBG+ZXfupx2RQFKg9wuGe/XaB1G6z4gXLIGSlvWJOhRGw0SLuyRPR2kxa+SgVC0m/kOMMh2r
sQjUiFW7L7VFuydPNd/dsZFOg1HjdvxF6lEx9NRP4okVtA0HcYem1iauX/Bxls5A3jYerLisu2W2
/QDg9D+oBh0MSEXQuCm3LxaSVeGb7ORWQ5/8ADna8NQ8KJSQRD1zGMttRaPsCdTKMJ2FYEiv7/9a
AGRmK03cIJWWIlkMDELEGD1wFDg4eCs7E0Xk6lRYAd2zTx21Rh9rcHjEC5bWEkb/SfpQTbYSn2RN
Y384Tuul75CUpcRTkeFh9fzomso3pIJ2YQvt2DWgqLiqQvnrCkCospa+x+JBZrxTVxZclI+JuoSV
A+YQ9BM//mVlouLRjanxYEnRG2npDhlRXYrsvAJN/Ei60E886pnX2n18IPTChYVlUoFG4I5xnbXJ
hjIXkBYuxaIhO6Ax+YWAJj7r+skp9mdb+RlzBNcSCZ88T88nspN736A0V8mW5Wh8M8nF+8A/vlji
IbTI6VXS6PPscq3Rlt0az6mpj+vzAxwrHtWe/+c6cdSD0leyW9CRzVp4mSybGaPmaHoYbkHA2+o1
bgq0bJhha4XfC64VvTeN+T/zIDJh6kX35Gd+o9gZVagwEjjG35BFP82FMuLNbi4QYnFuYo34qcRq
jXLEkqbmZdhEBNZFsjUmJxzPIsn+261H/PXm+PnN4R9UKieTroTNYOJIz199KE1jWB2XtfrQ42lw
pEJoUY5XpeDFnOGOX9sdNV9ATjbVvLjMawG1vISnwi7xieKLOsXTCIFckCXddSicxnMeqjVZe9cU
mjmhlRiD2FFEMz+112hpCzxJbBb95zT82K3p69malKLf6e1qUbkIv+z37yw7XG4WOG4rhWZ2D/c3
fNQ/2T++BicHzqjEzdwIujnRlX8poNwerEXSPBfL5WHxeHSh9eqgJn11XhiiY0hVixNu0LiN13Vd
RytXrPSidEebC9F1qJ+PiyXVoPoSSwsW6tMLtMS5MFFRdnuo4lAB59h/tXrS19Cc7aClNjIi2cBl
SX2Q2RVkPclf7y4Xa+pLXWGK2QiJD0Le6T7NB6dy16v+dWSalkmBZHybSUECZpVfd4KVDPzcerwY
nOPOfV/et0wLMROrmMmXD1fDCwcN/I0W75z86y6CR6V39IM3troU907Nzd4USD8lSPNmlOvPbS0H
ORK7UMmeTLAIRNfikfPX73FICVWMO4DfMfQLNoYYKWcK87+FOJofI1PliyqqjKtdndMogZzYlZp0
3bZgD+nG7gLhi6yty9BcIWY4vPBjVuekEueFvsEep3hFKAotSj46k+tt6/4KAm1OJBDDirZncQTi
gIk9htrnu9vLy1IhV7n1x5b4V+N0jNsfnzJ812jMXhpPAdiYWWKRIEanAa9nXzntDoI9G21JXLuf
IwVJsRRQ5QJg21SmJDwlo5HeMzf5eNnfRnBrYELoPTe3HtggM7GXxbStiRB+T81uItyyH4BSjCAQ
TCySTazjFKCuTRAdpXhy2zdKeoV3Scce3ObmvuBtMhT827h2PITqst/TGmKqys7yRTkeE7vaeAxn
MWtvAff+YrJ9NMXaOjWmXJ0d6o0VVYcZT1laYkALO0i8FljNAKRGUW/AJYKhxVTTrWPBhzMe24GM
4NKnd5b+SgAd/gRENehPJFkaKF97jx6J24RGY5CQsOnyAunHtuNjl8YCgZHfu7C8J7T2iAUqsrJw
Vf/WqxPck7c+oKOC4/7Wgo64kctD3wLiv3rMu+nT9GRc5oegLbpNCeITbsKPtlOjFtDI9obSyVgH
Uj/sS0l2Ip14Lc2ZV2e7cysUvrQco+ubsTLVPlXyf3kDBP2n3Phw7qNoHEqXNbqaDnGY7pPKSgLe
NIqaHQdlmbJgwe3T1jAYai2jtHLbvtzI3v7496teDf6TBcUZEmqN3ye90gwcygZx68XCEsI8Lwbh
0rDMoa/GxEXMwiQP2x0C+YLZXA3CnnxT3QX6+H0cvwSQwkZB6a5miUW8UOD6l4YBWaV6TXvXfKRJ
YGIilkfIfZ+6a9D4hcMnM9vKWr+3JaiwDc4ueG82/HG709nZiXnwWJ1NDEA/YYGdYP8bH0OCvhhQ
MIhJizBVMJLfb247vO43qzl5qCFfnXQCxaombayC0VotxMx4jXKhAAFvi8L+NHY28DeSNLNoO5o1
K9wa1FDLZmcZtjDz2HYqSYzhhhLCC2rPxI9kq3BJeu2mK0FCM0QGGnc4H4eiUmTazYsaEcWIFwRo
7tAmMAISpUo0V32IBJ4M0nfo84pX9zYX5h9PYJXO1LqwJph1nVqwIHSODIBNAZf128CDhxa3+ge5
GIoTmlBVXqo1I++kuGpbcDHcAVPkzRHpRmDipgFNsgCDN/R1zUuHm9uQrf8uiUO5ONV3g7uBrMjW
9mN+1SoHBYbuO6mmKtWYArqdbVqKwYJXlDSffOm0hl8ELDg7XVnEwUUIPaaJav4PGdGAeT+m0zfb
dHxc4h3kst/AHoKztYmemNoDYBn/MY2rBIlQRMRg5Whj49RD2GJ46Ojo6X4NjLVtfg9GZ5mVKgwI
yoVNSdXp0WSIEump2i5zeVRGEf7NwdzdDMTWT8aEo9SRwIFA+G1wmTbQC/MiHdI4a9sYYTs9WzWA
96L+4X05Py8CfTJMa0PQp/7bMI+3VfalzFIaMAwoSfKHLmgXnEodIFc+jPQ1RB6QcExniYcu8TdW
MFoFGlHFq3wttHZO/MhSjQ1rfJfJt3N623w5pyOmtgzxoTYYqKXk
`protect end_protected
