��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ��E�[2�����S�'��t�w�����b���"h����T�õ#����p`��0���8�V�b}��SV)ڿ�_a;�W�q�0�1s��e�v�0��*%G\|yN�@g)_��yt|̞Q���6���I���(��2$ںv͸8���{� gm�/2 ���郪�^�[&����a��o$nfXQ�0��.%����;լ����x�2g�`L3�NAgAL�����歲���!Q�Lr;����vr�V4���������l��=���n� �m\�
M��<�(�%�"�˰K�-��)��	�9�f�)!(Y��gLHt�V��}.5G��.+Y^Ju�t��1��I�+�b�IG�c��|��V""��v��UF��ڤ���� @������'.JG����B��9�I�Ȥ�s�����y|E�]N��=M	��ш���*��d�xz�
���c����m���,������$����%vĬ�?>��o���"�ZV(�8���)�@	��2-�5��O�)��_���cD� g�ͤ��x|��ލ�Y�jY��@j��S��5�;8\��OvK���5X�vIE��Аd��bQ��:������Dj��\.տT����Gb���Fx�m6�>�B(�����gU�$�d�u7�"�Q�蔨��?r����T�=0ɱ]��H��<�����xc��.f]�:��m��IӾ�BdW�cZe_�T�%��r��2l�*!�IOHc�8�!�H
�n�ѷ�oV�G�fx{��5l��d����BK�"l;+(z6�/���vm����*���%��:N���dq&4�5���o����o�:��8r��׬��������`[�y�)��S����/K��'V��\�N���~[N԰}?W�I�ңIxNm%��YT	��g�lʡ#&���nnv&~8=�ms
��V��a��V��"�G�,v��BƩ�o�j���c}�� �������d?��J��Ћ�����Z��6��ni�xi���CK��V�
F|�/;TX�g���c��N�� y�V����Rs�-��T�5�V�,Q�d����|��]���*o񐺁O�'�
�C�DF�f�\%&�kw�eER��F��r������ѹޮN��#0�~�b �l����k{'�gV����)z�r���IFPp�O(��D�T��o$G��0c��,;��u�R�R�<��]�sL�o�>=��!B��ݰ��kY�Sv���e@A{��P6�f��Ȏ�ý���&�6���eg@Y�C�:	���a��W*w=d����`%�}iO�)��<��~�������*?�=�V�.y�J��nк�m��jA<��d�uM�`��#4�����y�ڠ�L�#����gB÷��l��G�d���e�(n���1��v��-�m���3������o�jPU����y�`FbDz����H�� k?��N0?�H�{TKLU�#tb���nM55Ƌx� ��l���};N� �oC铩��LW)�ex�)RQ�[��3��.qA��
Zr1F��A��g���ҹ���������y�~\U�QT��}|���6X�&�+��d��;�	�+}����zP}<�]T�8l��){5�
�˄ڻ��5��g�L��@����,Zp�����F�8<1e�=O]�_�J�f��}��"�X�`�A~t2���^	��G���')����h��`���=r+{�K���e�±cH�1?�8�m�4��`���q�&�;*��Bb�zTSm����-t0h����q�=��̨���/fR��A�SUI���1�w����:��*Ÿ>���Se�;q�<�Y��b�z�&q��F'�D����r �33�R��&��_�j���� dro�  P��wC�~����Q)�BM����;�س��n>�s�B>&U%&8'��鳻o�wJh��X4iQ_�5ʰ��d��fO�΁�����GqY[|^����>�� � d����n�y^U��jW��U6_㹺�&M�tټ:�jKs~�N:Z��L
�3����/F;%7�)cʬ��=(�1#��ĭ���7��P6}8��/U>&������'J��N�ao�����zVgN!�ysW5}�$��]��O��h�nw�7�C�H����ܞMe1�zD`�Ix�}#�������y 0�AV��gT��\��v����N���;5�����X7E<	����"��G��}8e�|�P�0���"j�y�&I<����
aa#��.Eٝ�J��S�U�w�-.�� V�3>ё2/ 5��Վ4�Z��T'��/�g����a�Y��_�&�����p��l�����1�4$ �Q��H�,5K�[�$jq