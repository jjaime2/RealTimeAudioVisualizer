-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PnUa2Gva74CcjtwO/UU3X97nqlCLM6NeHveMhB6IyDeNvLw1ZvuoTaMTMvcMIpWsP+I2jevwRxRc
HhDwUNsgUfN8DtI21eLDLWsD7PxRsC+roD55VpMLJz5FvIhU6sxNSJ07h3qxh0KSoJEubFliSeIp
5q96eyTGp/CKV7O2BP1cijbxTXcLaKxMPxjeCxeorHvmKlV4rsbJHlrwiVNBAFtrQVtcZaNCfBd3
2XIH0lB/MhmKiWIpahcCLQdOMofcL5up0ph9zRFPIIP+Vp8vMo3bWgGtIGQnY/1yYjVg9Effgalc
gnh9rQqTDJqG5R9MNopvBiuWsT2HJO+XFEetVQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5536)
`protect data_block
LB42SGTqswGUY+h7TS/WCfzjN7N3S3kf1L5cmr2AZBwmpTepjfcqtXERZd8i9slbI+uYC55ADKWz
O9eSAcetd1kRiDSrzkuwHc2IIpTbp+aIVnnTozhCPKHnmNQ5NSDikDWGEkvqGVx3ErvPFZOltxjg
fK0bpDccK+wi93htArve0EYY4Aev8VQhOk40gm9RvVrd+fPD8nGsIbW6QdROisC330co0t25EWVt
gdvMh7A9Ams8XqWz4hjn81buQkiaLD49+CwBOXgy97+OzXTkwmuXlwTFzJsZdpgG6LBa/L04ddlf
0DcEbuvc7nqnhETDf2gqxdwFxMqiIpa5Kybp8hUuQ1G3oYwE1M9RQJl11kt1xwWtOEhx5jtEyClU
maKmkYyzgDHS8Saj+w1+NhXXoqLAvjBZBjll+vbWrPFog29n6wvZ1/LGifFgD185Zm0WHFZ8R2jV
cCPSFhRcLlX9S4LPJKsKroPLEowosZ6wmvF6spZp/rQtu1ijoSDlKnNur8Jr4zzg6FicDh5rO1JZ
T1vsX6mSa/u/K2SadAtuDSZfEXmEmpiMglUDAQEjd2YXd9Q+oN4nLKzpDY+TA1fmdIICkZYBY/Ut
iCooui1x2pdeyU4/P3URKUk6KK1EgDXjeAqbVsdBNHfJez53C+1Q/U72m0j/ZHlMkFv6SRkE4BVX
1ZgxI/xI5BEtJdLkJUAm/sTUH8gS+H8N7AKYSrZgVuVX3BGzIJnyjVN4ZU4cadUKatkhiUxyutgB
wL8BFLiwirF4VCfEU58nofWJNpKUF3BfhgYsgBq584g0AyqMJIKTesWQBnV9f2n+uU2rOpSuL/Nn
TVQi6dmiV4XvD+2Az6LuBRi1t9OlHFhRMZoaTdTsNlt7QH76lPb0ARJcJyv0b9rM6iCnKPMblczv
y4gukKa1CcWm/V5GhHMtYKsQV/pe/U29GuBCvUhoCsgKstUUFTv8/OthVbhO08DacuUaSMMctqoU
ME0BCCWgY9hizWnGAD/FdPHONbyTW3MqSjKC/0ZO4edakvYTK97kJgAAuzw00B1hRqEWc4ELtM/L
bgJ2gTvlZSzXtW3rGL83tH8Yrpxh4E8WMrLXWQNiz462ifGAOVChRBNlJntNJYq8tmpoG+Fwflha
zGPqRd3yBqWR4k+bJ7TpIymV5JBUS3xI2tT7EZCxSiIywH2ilpP3TjXBe9nafSgIaWqFnrtlaT1C
gtqnAzJmy3L8/QL3u3PfsDRx459YQXvpTjNtpa5+DJq812JeC9tvseO1z2y6AdX0KzueoEWU8FMx
PmgpRLKuA5POfPe7JaS09xVbE9ChATff/8oVUXqQpxavUjJ0f13BGsEuGmj13QtMaFXA0t6vh/V/
iLc603mkkszWlkdUnhnUrdFKR8K0pNgG7TCKqe3iD1Xgu62j8P1apciNCsraMWjI7zXzm5hbSQQO
HgaQxs5dfh5LykbaJSelsQXcO0vm3RNUjJRI+keop6TAPbRLYs74TZ7gAqOJAsDfkvWZ2vnv0TuN
Q/17RCxrJki5giOaEC47lOh43HGA6RRy8GwLbvS8wHk8yNvH4c0Mtc9jY1RVF+KMpWaTnJAxOPfw
eXTbC7dmhl5rQ+noKZh8UmoP/HqGV8QWgahJQcCRgkFIGkmEexPiRSMOnUlA7mtGQ3SFSDXgm4yL
SLciv3HEA743T40gpodfvP5p5h+auEMZkbWjdKD34JGuLEWoeeV4XfzAHmt46qwyoc2jtOrdgOcF
z5O8GrfQvyEVqfMHmUJMs5OP1G6I0Nb+MpOqueisbMZVqLnl9/zs8viIZOWlc2Pse2/mJTryglEN
vZ6/R3kOoiPNvjsUUY/BbD09lrFtB/6H6EqcL9kG4ujs01manx7fYZRKrPTRYh1m4r7lQCP8pfwa
8W4hGGPAaXckVOBA4Cs5kucht4mtwIFp1dQ9kKcdsFTvNu6H7WbvAcOxQVWsjeJS15uKjcVsSxGH
3LC73KQnZtVgs+r9VNPvrINkWSudgLyQKbL+4Q2qv65R9C8UkwKNfw5+XbDvQPNslz/sF3ZFxUCb
7+tY4k0Gstpg/zt4unFBfZPFpsQR4uvAlrbnZhzK2XG7pXRls2FQWWTX7hVLATilZDToYpAy4vv6
jGe04E0IOeJdcZow1CKGSIdamwvqDJYsBc6ArMi6LRfPa4qWrb8SdnhYEREd9T3/EMyBxxOukrV+
sQjLCZzFfFmczo+XpsD1MEan+w4AW4BV+Zw4InUSnNU4eYRNWfzQjcgC5C1eNRJEIg9AQ6+g6U7T
LuUzzn0wm6odoOfxBgM13G1Lr4Yc0jQLW98YUwWeTaz4vVz0eW0JPvhumSHfCLXzz7K8mqYKCmVA
+Bag4Yd6imZdzTzewtZwPhCaqYNOPrsq68/43Ljg+ftYZlDtXse8wG2TK5tJQJ+vFy6qH2hPvOLn
5xkkZgbHm4xdCpYIBKU0m/wyNO+XQvUZl2yPzaTbVylsupgDnhiqUtrJpk7q9FpUWMsKH1KESJPA
dpoQz2OH8uOhsh/GvAUDmFaSA8vRlL1m6IpHRgfvlPheONaxAXD4i1Bk3Y71uKTrBLYXWGitxZtJ
NCP7J9i25tX4yLVBQhq34yo07LtBzVi23eWAaVXsnd4W5Fcl1QcTEpObf7zlD6ot5Fws5ZERajnk
58ZlbSqD4qj7CPM7X1PKBKIooK1Eo89U9RxuakLBOgfJJ+MSni3BMj6wz/HJS17M0orkX04nf/3H
fj4ANcsf0O1WDj6HWLttIG0DvtJjhDisn1aSkIAyh+734NLpOnXDbJj48MQP4ZERL4Tf3x5YtsND
PVdZPMX1BtGCtgpxMYvmQcZZBv7LKTTACEcP07GqY74fRAIc91EnJiqFzh83/B0AybFxE3a4MFHx
E7iJ3xXWjxv6f36tPM9ebNEx4j/FXqPGRSHAZAfNcIrupke0Yuso70FStrl7QGOwGOPnK3GeQWxl
taU/O8JCWxlsEHTeh9bqc4vFROMIJkFpdyqT8VaeILCR9nilAQsJQAgQMGIxBJSz8djcDYIK0W9V
VM1ZOLiNvY2OLCZDVd0IOxE42+Wnv5k1K7mm9oG2jNfn2Naef1ql7/lc52Du2ARZF1V6Cp8w9FvH
efyYX4MdhF5hmVdHh4YatVFJ6rpfb6jTnJo7MGANEhsk8ylp+WkLQzrFuyDSTgO9xw24DOEYvbd1
2kVCYoeU2TS3p1omypi8uVWw+xw8KApPZP+0oi+hyTEUZfk2CEgGLnVnUyy3kf9Ii19Fh9Iuxq1t
5M8jbYR7IsYzOX5jHjPRvpjVOy4xS4h5Y1ItStCFq7Zw68ANnVlUqrYKLfiqksu3Lw0LN0ey8w26
gJ+QwlkxLM/a0+IiM+7teiOMc79S1izJ3RD/TMOwX4rpBuFCyxE/uKTnKkvMf6cWKRH2V+Gl5v0m
3/0uyauS2Bv2iTZnbE1SPYhb9pR1WFJcL3ovztYg+3VCaQchAFUnZwo+rLa/CArRiDVCIxJ3q4nO
8uwMk8PRUusaRWlULvCjRWGgwHVlCaRihDLmoyOsldsJacgxXoWTZdJf2o1CZIHSkMQhlrICx7dV
6D36dkXh7RMUGcYRKD2npf0kT1BeDfRBHvFU54PKBCC++W6MHRQe0hZMkJEB0sZ7WCP3VOI1Aqdc
bwl13abHeKFCbp/OaOw3KhFiU5trLbCNYAYIz83k+GvAqhE4+WPQuJ9bxbaTWEnjoTHElcV32f++
xVxxF/ilDW8T7BjQ+NFZ1RtXcxwW0mg9AHoTgvHJRA1ygKvpnBysVvkTLNVJGygOWEOhmDL8kJT5
MD+jHXAFtGOSxe0v8Uzl1nPReb2ray33ZwGui7FaE27GPJD4UFcRkopib+LL9ypEmt5Wdqh8H31Y
e01rXWXJIUq1aIU3NYMioo3b8FId/B7Rt2N1kNG2NO7GPvQbtQ1x2IhLHjj+WEzQszPR+mtLysvX
gq4thkjnfiX3UjkRzWo32jtFQAPUy0I5tXelAykgoCmBk7vgW666JOqg8Nrou+kVbYoAK/KI0ieE
aAOWTY44HhqJy1Bkrs58jVYRKh81/ZHNVNILpyH/cuLhntGvBA9JkkXJ8ahKT5UEuMa14/iMTWwi
3Zbvoi3+r4DsZTsPLAyv9iiD9/AOIm2MnaG5kissHL3U0jDstYlT2H0ufhASoY4TMYHC5JyApQ/6
usZg3hUXnL3yEVNFrJQJ3py46MWRt/7E8ZOdjPpYSEeovBtaiSwx7fYSNbuOrRmfNwDU/qxU0vzq
D96qEIGaO9DPq98ewpT8D/jSZCbZDFpn1nKYIro+xzPN8r4SEXEmXThc+v5MMlYTv+IkUTwhV+bt
VrkMJOgWB7Twvxt3xIMazROr2REzKeUmnLYRFNGOc6Ia9dNIt/wG0DKuO3k95CS6OofCeGBroSpN
S74MPHCfcz+cXJmGC8M76dG3g+TVNs31TTdn4uiFsx9uNvXUOHbAielhN2wQQVo2JnfLH27oW8XQ
uQB4AlNlsjqybWi3QorAJrpEqhDAIllp/RV+QrD2RlFrefMskLSVyfFHr4236wzvdYcba4KMyrhK
hrZyt+pXL+Yw3C9/sXaDNy0GI33fX0kQOH5HSVc/jivMH9hGNUThi85Ry7WNhzJOXcj+AeZDMUkg
ORzsei4/JiBVoR2IvzvWsC5x6Cx18WWddUVA/x/N+p0lXgeE407mEg5zFi7zpD3m2qKRdwQeq04I
EBqrh1vndLmlyp3O9ejD+1UdRxhvoixBCkqvO8LznjoKLxG9t3GD7HnJRFxI0j/5HowbyXuXbfqs
KBuinHP3ky9yIk+sVB3SE/25dfltQLKN/N9T1kmR3DdZHvPXOgTX9GNd/gYluhwnEe5r1HS+wO1r
6duFygUw8DnUfg/yJVNz/B74Y4NHh6loa5xEcsHFKlJXh1TdlxtRJm3AsgxGu0z22OadrhS/iKaj
eV2Ii/q2yujxdzK2D48x40xARsRfT7TCO/hj7HQVtm0/cEVXTd3Q0CzFWNa6fJ2mxW0NU0SogoOs
mgClHiOB679oO0dKSuWMejJfCkpFbTl+b2tk2i/E7Yn1wt5ODK/Z/5iQhEsJFWI0/jx4GkcVeSmA
kPCEwBY4jgte4xVFTTSZj0m5NoAS/i8oT6bEzSjkBfbuBTYmaiAVhjACYaJp24thyaFAE+EU36dZ
frpF5sRerYTYNdfUQQOkCfNskSCTuklASnSXeAMdKumchCzgmuJb7lBUuIOvwUQC5ESyUt+tzI5L
U0i76rLPQq40VrRs0uNHQRcS4tPALXp8QdkeTwedtK1yVhF9+qevanu0V74eDGknyPpY1Nrcuita
5jLUX/4L8M2OyIh6dPavGuH0QSA6Pu/xQG1Vhwhv9P5uIjDKm31a2Lqsm+HJ9teVsfb9o4N22xfv
g9E8GlH5frwVitG7CICnFm6rY6MeC7GUkPbJvt0EDzzLlDCglEAEdDSczOsTILc4f3V1JjWP7XFL
rQ88eRu5TUvJHL1a74UpGCwkiRAJeE4znAw6RoH3YkvAfDWYDquWCKzUGLrGAD1HN+dCkqZ6yH5G
evD30++rl4pZwo3SMMgGS5vodwineJZQn0elyOofY4ejhRRxOsKW3YIezchaEpTZZci3X8Yh9w+m
rAYNeng/zRCkp4zGJRsszrenbQbEHvfkT/dWWUorAue/bfAZTo0yfC1IJ3JH9+f5+kla2DHUjKyC
oK9lknIWhR+8iFfiu3/2OkWDP1+OEHF8EAWWZQQE3AyTJZe3hHtXQR5xtZFjrOt2CvXt6w3pkE8S
gkHczSAcoEq1lLSzBUAy1bimnNoXTU5JMsr3D0IlRJ3luM/mw0MJ2CJvbR6yYb9V2XvAFESDulhy
oBcybSiOfGl58dwxf3kq2QL0n123VOE3GvGu4/tq32deFQ7ZuJdfmAokwtJnV6H76z6EUhBvuvw4
ddv2LgF2PK8h5j/53SIEzRJfQwEalOrMn952rxi4OpZ6+bEyPWGYlhYdu6FYRn30FCKGtQdmoLSB
Dyxyl6MYC4M4RzdWYAQhwOARFr1nl1cnqlLb24IDgtTdFXkcgIFkXGmdAEOplriQMjv65C4JyBmQ
9QZLIa31C1P7ogm25zTir0MWq1mxHQgiWNaExmPTF/FHIl6kvw3swVrUQzcR3BhwE8/LeIK3qUU1
mCgtATCcVGc7SjIhHgmDXSUUGnRt+6Gi06fnFLxZ8czx8uRRmElMXHgS14CbtsCEnEFHkhEeS7Ex
cHqQ7E7CiE3v+My3eWS7QtfjjdbPuxjN9OhAy1HZBeBTZIGyJWhmhYMqDuNc1r0KTHD8yoq1QvWd
kmRQ7FF7/IQkUOhOcgnENAX4oOrF/1t3/hL8M+HHJgYEfnjulR28VBCnOKqXz86Y5KYzQsENd//T
gsKZ0hWIbPHcPs8McevvQ6HQYYt2orpHxQfDviZJ2HGKFHUc25Cwi0Rsb3pid04PdCcqlObA8Owr
82qnS9vocQ9UBiyvpzEEznLVgg9ow2wwrZKIHPPvl0ArOYUviRf9QomuH0w2rIX99Beu9l2J/AES
OIWShpS0oP33s2ZB/z18s0mfDatST9ZvlFaYxMXZ6n10vKxeuosp1wwN4DSFfIXTwwO099Aeimlo
uH0GoFZAgZpXZxpdui6u53dDBfc8prquaqHO2WTiX9gQWTCfFWsyfnZM0B4b8SzPxfzO0yaENkO5
w6oPP6iDPC8wqaBLBse+1rc0QzNsOcojGx5f+h7O1jTW7/e3Y2PUQNfHpjqQSNEZeh4zYm+Kg3Dy
pTArbGJ2t7xPeLJQfVy2cFt5m2ZIAZ6fQdGUqfugbHb3YcNfi0d6RshrQO91ZKX4atvSAgcHujKD
SpJa6dXFOXAA0eRV/cl9zRbu9ggwc1qTzGr0vojb/d+o6F9nLlGgjMpI4ASEpB3Wdskok2Scq0aq
sBn6+vNxVmXUXTxcbFbQw7D/vQPQQAJimSAhXqP7KpatdosAMjPlb4Dj2PlMZJc9yzQHhtwqnXpp
8fqwVFtOzUh8fjRIe8g30YLPClQSW5WLC7v9gsytkoumTA11Di0DfH7zk3ZBRUcpCxfvnGiaFjHa
bXOha1lMR5kdVAp+S0AjiKXHVoeUTxz22FHYBii+NQUDwLlJc+NXsO1Ytl+8WQ4XWzP61HD3VlRy
hn8HhvslrtWuR1hfrMpOwiKEZzJWiZVczGN/qqGvfDtU6Ka9ZAJz3bkUSfXioGnQCAzUpjzKqaQ/
g1e94r/InuBfWAVYPekYnf+sfXOhr76mSfpDvUD0rMHZMta0SktFdBUeiL66Nswz9EFoeDYOThqv
0bFe/n+wrthdYSfr08M6/f+YN9Fz7e9h8nMdMV9Sq1BFd94gjQsREsYepUOxPGHR6/WhFIPt/Z6T
tOMy/pok7Q==
`protect end_protected
