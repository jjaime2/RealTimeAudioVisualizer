��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊E����� ���u ���A�a�Neb�0���KQY���C���.gD,T"�=8"b"ݽ��	��oHՏ�����P;Nr�Ɏ��?���Bw�,~�VWj�:�rSU��47�mP����A��Gs���!+W��k�e.�U�>�>��T��|8ࢼtk�w��՘<��{ś,'B�$�O&�	1�Rh���K(xY�[+��ݠc���,�=�)ߝ��S��)�Y�1��L�����T�g���	k;�������X���Y��K ���*�M�Ƶ��,���Ų�P2ĽO��e���ʨ�]PXH��K�Ɲb�!���q�#�!ă�5a�D��;bI_�����d}F�t���c�6�o�>���V�$�K�M�Z;����e���@j�Mc,u�H-��3r5�n�U#�Ȉ:�a6��{^)_7!p\�i���J�����Lt��� y�ǿW���Ő�÷z��b�1�����Ĥ\$���'�ZbCjW*4�V~�}lE�@F��}�����O>�O�:��i�.�0�M.��kXo/q_،k�{B�Ή�$`�~	N9>8%�&{GaBA�(�,l|��ł��J˞�2]��T8If4+����7���kqj�Qî�X��8�ԕ��z�{��V�e^߈��׏t�AQ���^3�J&��b��Q1K\�ѡ�v�|=yf�/�)k:v�R����'��ך@s��M�}/��L�GDh,KdR��. bTm�e�7y��Z������h��&<(�U#���p�D'�����Z��\��� a�d-l+b�Z�Ί�8}/��*u�}��d4�X�����]�1`�j�qT�n����=�|�	�f���{ap�8�2�m�_%��ꔄh��c�UQA�Ž�Ȟr	+����J��nȆ��C\��P��aoVL�:!�5��e�{���L�/|�G )�ѳ�m�r�G0�|O~���@Gr��i00%�x��!��Vp)��+��%őD7�[�%"C��R�����璏R��_�Z��Xx��A��ӟ�W�������\��\�DA���!c#w���%�8�H���/��6
wz{�b��[�zvNT�7[��V�%�s�NީB�2�4�1
"�<(N���f����"��V�g�-Z1?�2`���,� J|�dK֖�y	�s�"��ܽ���#�����u5_�+�f���VJGw�ĭ�]�3`���"?�l����E��8S���=@~U
l`n�#��-��fv��H�~ha�@4��d$M�.t�
����Q��-�Yܳu��z���d���l��l���S w�΋K��R�eֲUO6�l�)$��D�v�	����3c0K������woY0��lKKz�,�)K�������χ��Q������FB}b�eSNR����Xӌ�}}(�Yle�P��O2��{�����S6�{2��ȫ�P!�'w��(��Ym��t��v���j���WT�_�b����5���̕>�hIe+�6�"�ʣY�5�,1�=3Xy�d�8�!i) �YӨ�[�4,�3���żtxR�+��t<㠩R$ƪ�A�B�~2����ͺ^ݜ_���`aa��N�L�ط�a�p|T��yIĺ����񎃅��'�m���O� {��H��:H+�X%n�rR9�;�i/�
�yE)kt���SR@��%� s;�Sw�/.�kC���h&�ǃ�([���Ȓ<�*�&q%�d�ż$�y��I����lХ6���f��4�1ଐ+� ���X>aUA�Gbum�Ba�GP��e�	�hR�q�SY趸+��8L��c���������d;��U�Z얩
Kq���6ge�I�m�Z�BWu�t�9�7�vZ����z`�O�3|NG��/��>ڀ�K�Ά�3�L��qc�ː��+W��#��U�B���O�$p���}��b�X�x�Z3^~��Ebd�W������_"p"������!a�����3N�K f�AZ㒿N) #�J��y �#~z>��P��aoI<�Q<���*rİU����Z��>&6�5Y����Ji���;d�j3빙L�P!B�Z�2���V���P�_�5<����}��g�GV^�b�S���
�$��TY��Lx ������P֫�1 �5ue�SE�betC�ª.�ⴵ͟�����v��J�����������뻣�dB�Id \����:��;4=��1�a���Zz�o;	��!o^�;�m/�_M�_M����Q�UM)��T�H^��	��"���S+O!��G�1-<�gP���2��9+ߟذ��uo�.����`\����C�1�|�YV]�?�j"�n�vvQ���-�W
KL_���޲@���sy�8��/cH܎;��)V�-�����W�����7�/G �f�-p�����"��I5���s_2�1��k�۞�~�[y����k' ��L\&^csA�~�R��ɝ��$b�l���/�|+�����l{��_)|�\��T17u�X�O�[5����%�1�� B����`�B�:�4��(O1ۍo('?�J:��M%0=��2yG']�5gȊ���T�=��t��7ZT�?��,��p[u�WZ��Zk��oe��tI}��+(+ڀϥAƶ���_q� ��}zx�o��Q��!�G�����T����joВDE��T��Ar���"$�Å���@�����=��	�L����/l��Q����bE��ܨ�+o_�9�v2�b��[��\+�Þ�|�@�#c�h
XB�;7������~��{ v%���*�弶��F�w_T�<�^��c����L��>��,;�DA���d)SW�M��B0�"~p�O�ZS�Ş�L,H� p��a��!�5���� �Q�(!�=S)p,>ۆ�&�:�L�h�.`Q����?_�}y�a���GDl`��hף���*5@PJ2��T��FtЋ}���]/VI��o6ƖS��es�ẅx�T��?�6�)�ͷ���v��E�w���ύsɊ�bUS�$Ҡ��E�?�=�V,�N@&��MF����q�Lo=g#�z��M` �)\�T�eJ���^��팁�Z�֛kȦ�ng"�S'�yTQ
�5�g�-Lb��H�fy� ����A���s���'uT�>E����\.�^U���H>�U�Je��%vx�P�1y�o���\)���=PcM�diw~�[?~\%EJ��(�ҙ��7h�"f�+H�>���j;��}��8 ���>㨛 �$�&/9?G��e��`�E��1D%��.�~L��������>�B��J���ړ����!8�t��̐	Ce����i��-FY�d<��H_���N���'�O�~/2B����=x�T�d' �=x͢�w5R$�]k1�yzq%6���T�y�ㇲ�W�oMZ��VU��и|駷��=���I�ړv
 A���T��ɸ\g�Q���[�`�),ɷ��v����"�{jҒشG;�8���5f5����E&B�s��7������Ax��R&Oހȩ�'`/v(;�_�HQ�&SO�_連���^�+Q�6X��0���E��<��$,���ީx'�&��P��IB���۰�Q���,��u�= I� �~[MH�3