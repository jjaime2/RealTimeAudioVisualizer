��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ���l�$�'�Z���u��E�a ��B'v/�γݩ%5=F�7z�N?ysV�k�b#!sI[-~�G�m��]v��G��&��qx���m/�H�w��V����f�Զ�vp��B��\6�Ads�-����jfc`�kQ:�k�ɭ�|��&Υ�B��n�R3l=���]�_���Ro���*s0��|Ft�m
D�e4,�t�N.��a�˽�T'�C<`�e����E(�!$r�)��}�����3j3Rċ����7@�(��zmt)�`��L���Ì���j�LWS�g�K=.����x���^~P�$�LOa�U��Ɛ�ZS�|�F���\��C�bS^�jDT���"PMwNA�5��6��*�ڤ0�*��b�6��Jx+��v1�B�b-��V�l=w$֭�?��j<�V:�>蚢@�t�
O�RXz�gk��J�e�p���Z�Ňf�dB���c���Nm�}}d���ҭеL:6�Y�9����tE��URUT��W�OD��=�e#�����&����v�3�e��G`��o����rB�~8+֓}����nTVj����E���|�	ھW�0�~魄��ߣ���k���Ujx7��`��	A���T��J��L����T�^'^9;��R_���3�v]��%N/�eBr���
u����ͷ1>�%�	���  &N< �X�<��.u�F
��O�헡�)�x���4ؿ��r=g��k��Tї��y���ҭ��/��u�r#~�X�]�w#;=��ְ���T�zc_g�@�۩m`w�Bŏ���ϝS&\td`u�����O���>�z��xf�:U�A}����U�D�c�����8�$=��,��mψE>��a�w�='�Zɿ�
�H�X唲g��fd,�� o���{&�K�d��| P3�hqko�R~�A�i`���d�4�d���o&o�˨�.�6�_������[Zz0�]@U�T�#M��ӽ��'�%�ܱy�_��^}e�
�:Or#��]=f�O,��9`�%ً@����m��T�fc��@}fA.��&�ؑ�]kid���ƟB�|ZĆ�8�Cx���A1Ő��K[lVl*�J�4�?) �˷�&����0����sm��r���.�4/�"&1�����霖�j��t��T8�ԹWn��ds^�҈�"�c�g�ic6�L�Pa'z�U�[ͭ���V��![���uG��I|��&b�fR� ���
��7���_2�i*G9�e���ؖ���;ȉ�a�j�~���
�@v��''d5�c�4��-���c8]ů⽕��G�	:\�\�p�%Y��eF�������%~ZF����F܀�����9Kv`(�>��I��p����8��4�=��]	�"�gPu��Yk���xQ|�7�p��@_v�$։=�v� i��Bm�u��=���2(r�M²����*MHa�v$,��T<$g&�,ᝈ�  ��(��a+��2�놖.w\q���s��g�o�?�˟k$f�Y�#�N���4���e�{�>��c�Se���~.�1��:~�G��]Q�O)_u��K��D�?�j"��?:�xKL�.��@�?kP�Tca�I���G��T{G�,8~s[}�AfW
ڳ�|w�8b���Z�;������	�uw�s�v C[x+�weMVh�z�Y�!Bjj~�w�Jڌ�u\���֎b���`ۚ(B�QH�Bsq1[N bBK�׆.�3�Z����@�IL�U�@�3����X�_��5��h��_	��0���b{s�f���-�CRH>�	D���Q
JVf����s
9U(�^/@��U�e�Ǡ�%�����!&h��j�¨ߓ�<�' lE]0���I��=���*�\&v�M�Z�ؒ�|��U=+���.2`�8�{q�~�d��ѥ�IuĊ��+^\��L��O�m�p
��/��m���c�Xnu����f�	s��!Y���`FR�����e=���`"�s8�.'=���v}��Fy���לI�J���,S�"�ڢ�|����J���*�ǐ���ϮjT�cd�	�z�SP������ɌgBĆc%Fs�Rv$�nΑ��%{5�Lq_f���%�����'z�I��ņ���"�_�į_O���	�-.�.�Yb��1��_�[S&��io�z<�륛���)!��ȍB��b�4�-05�U�z�f6��ۆ�'�6�)/k�UN�2&#�l�w��!��� �W13Ɍ6obPT���g��ُo�c)hY	k�3B��w�ԁr����v�	�
��rpN��Z��K��F�T�����¸��'Sr��>���v`gl���{b��&M����Ň��Y���O{�ad��>$7\�R�M�8	Rcr�\y�\�6z�~��:�9��a�X����xOп�����S���1CE��0��@*p�h���i����J��?�6@��~UD���� �~9ok��5�O�d�r�rً�@� u����@q����~��
�ec�"%Od�+P%��o���=��1�������x�{L���T<{2˒�����ǵ��CІ�*q�z�i(G�FЦ�~���q�WX�\�q�������*։�=V3�p�i)_���x�2%p�W7�
�`�������M�@���G�����*/R �j�(TE��1	��o���Y���-����)z�!V(A�����3��8��?*]�Z������q���m��=�|d�sR��j� ��=�Lis1������]a�j�*3�����Upg���St��5����U�C3\�#/k:�$@�[q�G�ucLuE\��s=M�}�u�M͡z�Z�B���m��M3'VZ������@=_`x ���h���o���&uNQ˾�<�(�V$�U~��2��G�U�D:k�1��*8N;U��hެ�/�$6|��lF ���Gid	$t_,U�IP���\�[iRˊ[��B�w�_���t����W��J՝�x��Z	yRx��~��Sɗ�f|�!d���Uu�A-���|�E�5��~͎��>_�]]�	��ě[�K���x�̹Y���,.�kh�k���v�2���Eed�C�]��������{Nq��+1
���N)�_�����X��`j}-@��-����%�*v�r%4	#����`n��md66\ ��y�7=E Y���un��0ؘ��F��_g����p�����������IZ7�8sIe�����5�a�l�h�[0��pt	�S� ؚ��<:�\� �m��WX#�7��!��mY=t�h���-��ɍg�;�*|�ZG��.P��78�]�e�I>�y�I�,��T�̎ː��+c��wM������!{>��E�=5�~/!,z<V�22�*��;�6�ڟ�Q���<sX�"�p@B��3E����>�=#�w�Yoj஭9s"�&�3:gŴY@��[}�z��Y�lأZi�f�? n�7r���<[!]Ȱ;H6>a�لA��tv�'�`Py�ms��
�F@#3�N���Jo�D\	։f���v��òA���Xl�h���Y�ڂo:�ե���-�}G��ˤ]�_�S(���L!���������o����"z���e���U@�9e��Wn�w�XW���ǟ���2���(�)�`�v��k�^����������]�+��`��Et�,4�LE��e7̎"R�ʲ}
ȾsqI�e|7�Wi�'� �v+�l��?:����(�u�`֒G��'�^��l�^����m���� �A�.�ۥ!lH�1ǕW*����� uj�X@f�~�K[a3�*�33�R7�>cj�����R�қ�j�N\CA��-qzC8����p�V�nT��t�����������0NMm�|���C�h�ۍ�&����R������&͗e�ҏ�od�4����극_\�a��zD��pΠ�& �|�h��\�wGJ�����/��6����t�Cz��)~@i,��߼�r�	�P�@�ۛ�\��c]
t�9��o���Xz���E��wRW���T{$�*zC-�O�|�ƉTJ6Jڬn�������5��U֔�P��� Q��}��b�m�P�};����Ƚ�dñ!9b��+����j�Y��^��|e�-�Ǟ+�l3��'zɿ U�|V C��sY���ʕ��!��%�}��!�	��o�����f�ׂd@P�Io}�2)Z	˄B=���J����1p�g��ʧ�ï'����]��E�?Z8E:Z�ݢ�P)M9̝�xV�1�m���'�T�_hN�xI'E���	5!Ѐ��B~u%�ؤ���o�ػ��ׅ0"�N,|Gc"X�� ��n5E-��*|ņ�	G��ek��q��k9\R��~��.�������:=�y�Y��1I�CIULq6�z���:%AW;�7q���T'�%�<d'r�{��6�:��{�ۉ�;h��VL0*1ݗ����Qb��x�;b7�%%t�g��l~ㇳ:E4�3�l��H	��cqm{��;�'=��SG^�&�l��@1 ��V�����F��>	��2=��{������5�H�)�\��Tz!�B���x	��k��esްL�z�|M�иn������pU c�I�z�u�+3�l��fY�.�H}`^4���H{��gT#��S�(JBQ�E��C���4�UU�d^k!���lݲ�a%��7Qaغ8a.-m��ܫ�BLF��
t��q�j��s(�!D��1a��4��SL����,:�E�pدp	�q�1oH��ɪۺk[6K���&��^�NO��Jp}���U���CJm���O$͠ϋ#��xI�?����D���ͅ�ܢK-��6; fha抿i1o�s,��#0P �EOA�aG'����+�d����f�.�"Ap�+jDRF�[�)R�("�;��M"כƱ^�N.�E0]��6�k�3v�ƭr�o�w�ȿ�x �A���F �e�c
�j�����4�&����%HkE��a�:7?�w�6�Y�m�X8��SR�F��tԟ����j�A@AJX{�� RY��-���o�`L�1ܔ�����T�ӣ��;��� �E�w(}
����	PG���Z~w~0��ֳ�W�:��c]6��'��HL��n�����Ic��Y��8�y�љ\)��y�cnTٵ��0��p_�JTy�������à�iX{H��~�Q7z_�!ݮ�z���~��+ToW���g!L0S�
�Y���8�y����9ӝ�#*�ĝ��,�#�T�@�V�W���R�~2�k��	��踔��a��tԥ�/f�lY��Վ
�s���K^fϩ^���d���i`�w�hd�j�ԿҥWv�׽�GlM�P��2��v��?���]M�Q��T���kl3��vTď`�E�DU��DLn��QUGE�����
$�M˂�3V�r����Bn�O��Q��e�6�k�k��y&~�]<��X��K��^u%c�q�ˢ�M��ץ�u�^�yu5 �R��.�"��I��kd���cW��옣rN��{QJ�f���K$���|棰��6���)A�f�0j���צX�J���.n��Q�8T�M����$>�<(�6~>di�]e�u��{1�����
b�[�����`d��gPe �V���x��37�mB�܎J;�ڴSj u��Y}=�v 3"\�*��%���#�-旛��)7�j��i1��m0�~�sOP��7&�	�%ۂ�$T��Gl�7xӕ��@SD7�tq�
��n�p3C}m���j� b5'ȴ,O���)Xq�-��M9��}U��f㱇���\�t&�	;���Q�zK�{���o
!��\��>�6�Y4KpA>����ܢ�7�ϰ�����نW��<lb�Յ����0X�01Pu�R�����qO��k����~1=�C��D�Qe?���	SDs��-��SF����E��	��s�t)�X��8ŭ�yS<砷���"���3|Lw�\�0�̑˶N��6�ߺ\�ǂb��~{�ا��+��:U7��ۂ�<i��R�1Q�Wզ�,J1���
-�l����L�g�8^֞i�?
'8�7�C�O8���L�&'<N!k�=OзE��,3�8�N����qˎ�xx;��V�.�C�g����W��eȐ۩*�Z��CKk#=cA�S��<�0mE�#�E���(�����."�@�X^<�#��/��߅�=�j;���^�;nЇ:\�����k=vf߮86�9+�=��;toK�޳w$�j4\�Lŝ��t*6}~�1�8����I8��p�j�r�ك�䌚?�e-���o�t�}d�O3W��KY1�HOc�]��x�(@淅��'PW;��LV��R��)n�:j�S�Xmy��m6�M���q5$������\8�ў������#��A��4�q�$k�h�����ba��^it^Ktv���Ƀc��o��1�a^(��h��r�/���ㅃG��h3��FB��ޕ��S��)#z#�qT�&V��ĉU�(�gd~r��XK��Ih
D������^x��#>�q�	���kb�}���J,��͏$\��TZ��b�9������ı1h����PZ�#��ԘF�-�4�	�W7��T�uO��'�U��nQ�Eb���@t�|u���G���1��,�<�U$��t4!E9*�0��<�%����D2����Z�R��Wn��_�DrÖ�����[��{,���WXD��}x��!��\S0�����߂>�	�k��hBLG�?`�K�x%������\�	��}f�<�/����:������JS�+�;�V�''��vb��|�]Q���8�<�j6�����0��(�2��Z�4�h&|`�YQE� �JR�{��F��בBn�_���,��=DD.�:�4N�h�����'΋l��d�z���|�\��Bdy{^ldzM8 �m�-=��tM�ť�`���ՠFw�$���Baq�vw���|�9��%!(�:XU��2_�rP���5����)�
ˋh)=͑2.ϟD!�bj���Q���7s��$ffA�g���4�}�x�g�j|��.�� ���X�ccP71Τ� ;X׊1>S�Xua@�!�v;�߷	;��ѽ�=zJ����9hX�9 �$ʇ߉/�]���R���	+vAO^��O�8(}`��voQ��Bn.H0�ߤ�3�e��g�-$V!��ȹØ�E���@&W�Glp�Ju�vr\�$C���#>& �*3`{����:����CE��E�S�F�
�LU�ڄ��,��~i� mp�Ϳ!�
��� �_���l�@����M���:u��:гB��m	�G�΢��ڜaq�wu˛��;-��_�rp9d:.s���_�k>����(]n�jy�0P���w�]}C|�<���<Ռ"P�������]ɪ��{f�yT�3	����|`{�qMlo�Av�H~�c�8d�hQ��:y/^1C6���)�^+FOj��	o_�>���(yģ&_��!�-:����$P����K���K�#�mR���
B�h��B����b`38�m�1�Ǩ��O�Imu��H��RB�L��ʹY���u��d^�B9���jI�+a�&��T;��P;	5&L#ڲ��{�~V�Gc�V v$ȥ���P�^�4&�յ6�y��z�o�6j��k���isL�T�G�;l��T5����3Ϣ��n.g���=W�g$�HQ��!j$�͈��ʻǨ:2��5֔\D���&l�������!ĭ��+ U�6��Haj�T9l՛� ӱf�d�4EQ�_�J��"�0�n���b�zi� j��&�p.hݚ�'	��l="��h���a�%=W�L��j𧃼�Ť瘔�J�]�e<���V���t^��qB�L*��#�,��?-�z�
�Or}7�96Uy�u�[t���M�eJ�ـ���iw�f�14��/
����rX�����D��r��w���m&]�W,8nf�(<a?�靰�I��B��>�ʾֻ#6�hLM��}1zU}��>�wg�m*N9�(�˓*��]��7�kb:Ӽ:��JB*!�<�!,�{���#�ۿ�]0�NmQ�pF�ԓ��5�~�-�Oo���*䙂����Sȁ2���}�z�z禎L)�h�H��?o�4yZ9�'ߣ[-+csY��\ǉ/[���Dn$O�nY"\�↮G0�/���'Ms�Vʰ����P9��qٛ�eih���u���ͬ@�6�gw&��'L��(�,�j.c�>���s�]h�Tƙd�d�
��Y�uu��ȹj[�J��T�+X��_�F菁q+7�+��a��^�0wX��L�|%^�ÐO�Ԗ �����dnkG��8��Y]���b����o݆�yб�Y$;�s�[�ّ��t��z,h�t��?ZA]�I#d�5}K��z�F)Q��>o��5�
r�m̄����٢Ю���f����x(�u�m��[��7.�Nt�����Rb}M���b��� �Z���y}&HC��Q�x)Z�(�l_�3l���#��Ш9-��yx	�<@� ���O I~^��C�zc�2���bN!!0������
�Pt�G;��2�D��A��v�5����,r]r|��<�]���J�nF����ԉ��#]�'�p���Z�lIX�Yk���zo,��熘LOu�Uc8W|]Z�H~�yD1Z1~��°K�\l��z���Ͼ�1�f���\���=l^8���?�mn�tD_�����m0��1�F(\P��B����&9���h�+��Fg'��cn�!��)R�KT�L l)+LU���T5=��J�$�rښ7[Įd)'�[S77�8kɕ��.2bh�G �t]�K�:�O�Z�1�k��� @�!���.�i#�A�H��2��d}������2�{r��i� ��1�E�"��u�@I�-��Y��;���Un�-<�Y��`l�i���ċ*x�a`�zތ�"N��MJ�l��o���&`Ň�2t������*�*)]�D���o��{�2a��Qsu���U-�^�����#��c�I����[-\�� ���"J+r�`>uFt'���X�VZF_��Vc�:����A�Six��E�-������܊\�ρ���p��Sd�x�q�����:6��I��״M�1%�8�%867CKq��Λ��ns�ʎ���a�7��V�ʰ���Iw���J�,E��@�%	Y�)�`V�Qt���)�C��{ �މB����B+jM0Z�/�Q�m ]6��J����K����f_�h�Vo7lv[V,ƍ��������K�
�H��E�+Ʈ3�S�J�r���! vxƚ���v-��'�Hm��),�U�*�7&�	
�Ƥ������ĩ������k���R�;��>�*CM���5�Ï�" �5�	]t�Π�v��=$bv�&�[��5]�R;k���c�H����bΊ���&��<���ƮW�N����!�/�w"ٖ��t{Ha=�@��c1Nsh��}J֫q�a�n���	�^C����cF��i�+���~�� 5��r���������<�G��[�*�ڼ�Jٹ���E87&HV8��H)�OtL��Ɍ7&��Ye+%���Ո�����X<����Z�Gb���%�8��bY�:f̡��Q�K�(0�8��V΅Z���#}�z�*����P�(�6d��m\��i�m�Rl���s�>�C �̋�N�u��f\��v��1BOc��4�\���
.?��4��ا��hQ�������C��Be�}b�gW�ʧ�z��v�Un��:��aw�x$$+'Ȗ�)��/���136�+x��7w��7n.;,#<O(|�q�\�TNHC֪�tv�M�J����貥��0�O�ja�TsoV
iR��5��~�nc۽�%h0���'t��Ձ���J�"�(Z��<v]�tٸ0P;����A�(È�C�� R�
c���܍O��%l���`r$�A��
�B�c�37��J�$��E������(��a&�T��ֹ���3�a�HD�M�@D������0Z̗_+n����6.�����<��pПs��0Q���5�;����nL�).�&z����+_�6���<:��.�y�D���NOlIW3W8utnဵ��^"�j�Y�s��[��I��i	��%�Æu�1R��(g�o�_r8b8r�Yy;#	Yk�-ϳ�g�u8��������k�'�J�ˑ��V��n�y�_Ge�K{���*�Vs�y�-r�hg9�ٓ��o���ñ�C�r�#x֢���
xI�9�3�t{���s�5d#�	B���5��PjJt�� fvd� ��?�f:��"�nŌO�|S�x���J ���
���zߪE��KS�W��o��RC{�]��da"���g���$����H����Ȍʯ�"���
ׅ��q@��W��]��ʘ5����}������QN�9��$� zQ���҉�:Y?&�K,���=�1�ʣͽ���)�7�x��9"�	��O=��J3�����_Z�- �5�R�Ղ
Q�DG��T�^8.Ǘ@^�O�O�VRd	�����v�S�M<���-�U�v:�̢Z�U�^���u�a���	���[�\�6�s�^��҅�8� �d�3������@����3)���F^On�1���-��2a���۞�tBA$�R�jUKts�֑��{��
�3�B�a���KAv�}*��r)����ش\d/�Gڢر/&2rӉ_W辍�d-x9�9J����X��p���d�D޾��h�{���"�-z��q�b@��z-s�Q��W2�(�W�$��Z�{󶤹��{�f�ĄB�����s���L{��q".6��SI�yI�e{'�D�İ��J�6�Z?��ČiV�p��ůiey R�}�y?΃b�ڌ8ݘ$>�Cp�%�<`�\M[���`]z�5���2�F�p�qk�<�i��&��|�p�좚�¡[�2�[��E#W���9���f,4/Ȟ�f�Op���~�#�*��P��u�з�I�9�m
�[s�� ��f.ߪ왇��6�	!3����4jޭ!s���
�|�/vcuG�]��}{�K�YDI�E�(�5^Z�WJkߡ33��G6�LS�����L��_��ݳ�+%��'�J�vtU�5f���E��@jA���#����u��מ���#�5'��z�ŷ�[�'ʞk���DU����	П9/�ͥX�\�ο4oy�l���#c� I?���4~�$��&I�]0,�o���<�<Z�j`T�?]��W&��Gie��g��q��-Ǝ�<�Ǿ�/T�>K�V�����(R�rw�7�ͯ����*O+��FT�킓e'����
������g��،���0��V�R�Z�6�|�M
�5n�3ٞ1R���p�6�����k���@(>[$2��_<w����t�l�� �F���H�!A��hwz�I����"�hUl)ˋ�m�)������,�g�s�O�:6k�u�p�V�Ezg�b෧����P��dM-6��He�_�a�Q�"�M���'���% ֟�G����%]ߞ���\�H�zY4�S��S��D>Y]���~��ӹo�����a�t�ݥ�n�}�a[�&}����{�-UI�B`H�U��
`iy�$���!p.�ͤ���1S��P~\m���
8 �(�m�zs�+�r.~B()*�+��ړ�����#[p(��IT������"̪fk�8�w��g�z��_��w�
E(W�"�́O�	��^���5�����	���ַb�n�q��������@!v��A�6��lo.V[
��6��@���1�^}bVE*�!l
�3Eհg񔗊\}�dEz�����K��9L}�ɦy��G���h�g'`�k��h��a5�j!Wݰ��JE����۫�R�/a���邈��Y��nH²}���2�h=V��_o(��wn#��1D㱜�a�r-f_?�6{<��55�������2u����WU��Oe�JKjt��%��g(���'[��4`����������@�����Ο���/�LMds��p��n���٤$�Q��;=�>�
���C	�i�,�� A�ش�!�Z�g�����ͅ���R�H+:-��d���v��0.c�[���~��C����EY��	Ĭ�_�D횻�1�A�Q�*C)�F���Dk�0��z�I��ۜ`kD5j+�{J�Z_*	�ӯ)H?����6(�W=Y�f�$)��;�p�+Á�"�M7�����K�t����x?.�����W�ka����r�[��VS����p�tɺ5�%��m��N/���ָ�xU`��l ����C_ ^�:w	%���/�w]o����^���`�!�+�Z�Ī)��Е���q���W6T�����,��Bsco��;�%�;��]��T�Pb�j;v��|�M���:=q�2��'��A?wr����R����Ϝow1����:�Jke��u%�E�ڹ53�¬�� O�v�b�q��¸1ĦO:(�(�d)�M�z!W4�"О���5!}�]'GpT۝(���\QV�����,0KÃ�]�[�2�ue���-�vE�\�h�<w���ڟʪ�l����䣚����DI4o��|'8�<��<��,ܘ��׋�\�/���o6 !T�yec٤Ti.�v#�l[��{O>"|����8O*3X=jN�/ �S�m�u��ݰ$�?�
�1�K@X9��4����z�ۋ'�^2Bq��\�'����N@�ͣ=yt�ﶘ� �a/�M�Y�P��ڞy����Zn:%hcGs �S���6��.VJ�ix���u4�-I�����..$Am�x��������\�V �yw�'�oQ���`�E�[���r���<��͑��
W~��J�-*栖c������ �@��Er��W��w���	}��Z�ב;�p�\���r���`��kCW;�&P�G1%<NM�#�#��=<��qzќ�y���W	���|�c�m���ynQ�	~ܤ|�\f��}zy�_:��
��4�x^e���'��;ȕ#�^5�E�u�W��.��P��i(a�b+02��N�V��VlJwo��c���td��5QÂ��`%�가�����w~�W��}(��4�	;.��B%��l!Y�T]�����	��-�-?�G�'�4�c��ܖb��t�r��3��K_#q[ɰR�b�1�s�<h ��C����K�Ad��r8� �E�����Je���s�X{�eE7?������p��L�`8�%A���T�>�ʚ1
�� ]i����
{NX��IX,�ۺ�@l�"o�_�{S7�fٕ2���A�����S� �m�i�e�Q���] Luic��U����:e���v8`0Lp+�՘���~~t4��n��G����B%�����/�\�CCm+�6,��)'��}����]�"8p�)z��3L���aش>u"}��O�A.�>�r��L Ѝ��������U1�mk�9_[�}��IӹÄK��aM��(�Z�)�S&�5�N̳���� ~:��9X����?���H��r�,?�{��>���y"�^����.�h�������� 9,m�d�{gw��>��`��.��R�[��\Y��Z��=�n{�ߝ�`��~����Q�s��b��9��J^��r�����b��Y Z`�6?�_ڄ�bO*�^�$����Q�����Z��
i�j|E�R��|R�GI��UDK7�m�r�� �AaכwZeo���#8�6�O�g��`5����L@��D�!��-ï��k;�O'3�Jܕ꺚/�6Y�ѲF�/� �{�D���!F"�GR^�l�bo�my�+���~�D�����F!��	����R�p�j;eۦ΋��՛_&/�����w��
�9�m����/W��K�*b�	+?�[�,�k���Mi륩�Q,9Q����ڵM�v�kx�"\5�T�W�/p��cH���A���}�V�Xn��XMJ�ȷ(P���ŠO���W7=#I����X*���Vj��y�اDZ��+���+��j�ݱ�r<F&�t3p;��_X �:�BW�[!�b��4
[]��j�e�T�ck}I���S���"xL-�C�x��V�ETD�
�n���8����^�45<1����vVW���U���ZKs&2��fb���+�l�=��wU:(�՜���P�1ZW��d���2	�0j�p��e��Ժ� :�4S^�U�اe]�Z��@���$[ȹ�ڜh ��Q�D�h��[�R���Ȳ�V+�/H��9��z�+|Щ&5�F��X���k�첖��]�Ĭh��捥�@�F�'�f#�o��$���Lt0/3ikK�CN`!��C���Y_O2CW�K��Į�C�Ղ}ޟO1zR�䄧��f�!y�C> �2�<?��y��n����"GP�����y�&�w<�B:RH��1���掚0%�1�; ���sLm+2E�0�ɒ	k$�� �M�Sf^�Y3I���k�[�`F��"���aZ�ߟ�E������0���Lѝ��<�#+�TV�+�'�Th�e��3���!��i~=%�jX����D`
���>	���I�F��}ԛHS>"T�j-1��S�Ɔ��h ������@����ݪz�6K�\�k�k���S�/��c���:& f�'�����IM\�In�.�D3��,�x\�g�-˓[H�՗�j�:�E˷Q�B�h�n�N��H���1Νy��,b��xF7ut���6� �F�<
hГ�0P����	��gA���}����*�+~���l��z7�U�7l7��߬�x=X1���6��H��8d�k����V��z~�j����5�����EM;RT�?ʘs=�h
��^)Er�pg�{�����ڻ�
	��ݔ�^;�Vl})	�cx�Z��Ĥ�Y��ի�z�ڞ�):>�:8�-�TӚl~��'�>�1��삶�S#_��a�r5�7���2R7H��8[&Ӹ64�p�}}�{�T��IPn���?"�U5�,��&�W~j���}+�ڇ�{�HR�}�
�Sa ~a������Q�6�ɾ�Xm{�x�7��mŘ0��fz��$q�.�8���y�\���;���s�U�+E4`��\5�o�3�~��f�H9���y����w�6�o�Y4�h�����i�u:}��c���� g�i��*h	eկCFMf��D(_V��Ӓ����n3���xc��SE�YO��O���*L
��_&h�(���~v��E;����E5\,�"����[�	[Zg�R&M��׭	D�Y2cCj����Y�ꇚ�{%ʉ�k�,k�������,��
�U��m ��4�����u�;�.	�Fu�����h�H/��G����b��x����$g"V�M�Sj�E$ԍ}U�=��)��9Q틠y=:���̢�0C^(����A��0��B�#PZ�&��x��ȧk�չD�:%���V���9V/-��+�V]���rf�}E9���/���k�(yn>�L7������hFD�S�:O�f��A��b�K��aq	�jpn�b'�5���S������tn�1�ڹF�-jF�njc`�!��G��݂�K�ry��]7&x��2�s-��G����a�'[�/�ߨ��ѧ2%H���(�=��Y6�mˍ��	�!�\`&�E4�gt%��� ި6b�˨��״�^$6��c�38�D���8�1��p�P��C;�w~�&d�zmo���,n��],`g]˖8D9�0Ƚ�m� :7�Z�5����U\�i�$�׮$׵.��ғbu�d��1E��[����S��x*7��
��01�i��Aþ�ԕ�l��6�i���6$R�D�ʲN�Ȑ�d�~Z� ��]�~l
��5���3��?�QLB�-��y��v�5V��1�n�sTf���4�j��h3�����֒�E�R�ؚ,�%�IQU^����<�EM����Zv�7�R����wn�_��ɹ�30� z��l4��G��ઑ�=F��bfD#.����)9֢��&��I��x�g�U ?��R��]5αa)D�ӌ�H�B�K���T�#aQ�]�L�EP�A��lsE�(�j��oA�G�˔�S��sb�]�$_`W�=����5�Ԧ��:�F\J�]�g|�x݃P�}���Qk+�d1e��ׇ+��-��������9L��������ƤJ��(��`Z�4���@��cRh��i��d�U�l��6��� ���D����h�x��t������'�z�D�nF�KXrJ[}��.ڞ �ţ�<�a��r��Ԗ��:����%+�.��G�/�*����S+B�tXi4u���njK@ѽ��N3�䵺���PH�tڙ1Ǥ�U���x�R���-�e;0��ow²���8�"?Mxg��`��Y�jѓ|�iG�t²�\3�F�1'��?�5v`�"x
q(w��.TiȌ�����9흴	.y@8t�!��V\��SKc`w��B���]�;Һ*�Y�И�;$pl0:�!�
(Aq#b
�w9⊏�6���>�!h�T��)���t;���a����g��7Z�m]c�&@ՋW����"�z��#�`�Mۛ٪�l�����^��q��oqwN������屰���>,:=��k�̎!�I�edF�����j�7�]�d��#�/K�C���=��[��B: �mw����`#���b��k���
 �J��(�QO&Jz�#�01��	Z��Q3�,�j
l����H�+1|/�(����ݖq>c;}t ��O>x��
C��l7�R��C����p?��ߒ�bX� E�����+�N9�-y�W�0e�۶�Vd&��+{�b�i��D%)��^�-��r���٬��H�Z(��7M~��gc����J�i��C�W�3X�t��y���9��-�V_�� L*�X����q}��r���3�Ω}KI��}�V�U��h�u��c1/��e���{��95�+@����#f��v��K|s=�a����a��W�
1�Ns�.��a�C��~u�~�BKy���BU��"�磎�*B���T��Bʡs^`��q�R>�*z!:��<����^P!�Bj��:��s���9Ǻ�uG���t}z��7����{��	9��}���9ė��%_6��	�Pײ{��k���5��{}Z:�~�#l�!��Cy2'�[����:���k�|2��d��7��N��hb�c;�a���+>"m>�l��%� '�y�Jtu���~�����x�� �d�d��Z���ȗE�J��>��Eqon��±F�-�c1����vk��&4X������η����Yc�"��A#���m}�NG.Ʊ�1��!�� ��>�j=�n�ܙ�H�2��'���5^0c��Ҁ�xm��"X�5ƿk%O�bM'�4B7'�-.��ۘ��ů��D�����}�cZrʑ�&�P:���/�����z�T] ��I9��z�o��u7�i�d6SD�?FI��8�I�����,��U�;��Ї�ni���R�~��&}X��\/%��+pL?.N�m4&5��9a�s��Ǆԩ��R���1Y͗��Ч�"���@�e��N�6��|2�z��0�et��M��Jw��������UV���}�o�����b���"~+Y��va�1�S����N]ٱ����O�"5�r<�M%{MtR0 ������ BS4��Gװ�^H���;S�+	�k�����b���8\,�yǤ�%i<��Y��1*R3��K(��ȣ�.X��n�]D����o<�d�ȿ I�4��k_��	e�@������{Ϧ���y*� �CObTqu6�oS�o�.��fܴ�O,��&�&S$X��+�@Q��4/e]�r}�D�����>OF� �te]3 ㊦8D�_��tw���|&��0�L<L��y%�5�h慀W(�6�tp�M�$p^�H�8��i�	�>#���h�,�E�����<�\���DF�+y��잮j���8�Nf��/��+ge�q�S���N���!.֥�㸡��->�l�o���Λ���u��j7ϊi�;2f^��3���@z}2 �*���B;)�0��k�E����&E���s��GCG��d�{�g���M�6:>�{j|�¿����
jhT^��]��
֯6�A&R�\��U�B� 1��ҀS�7��KH߅څ!�������GW��ځ
�f�L_"s�����:������k9��H_��ʐ�B���d�g=�J!��QO��|2'� �P��7����g�3��'ڥ�l΂5��=,z7�.r9�cGz�&��  ���SS�ȮM�4��ּ��dᩲX���7Z$~[UV�{�F�ٲt��/����9�z{��|ٖ�%jW�=�p���M�ʚ�(�v�����+���c�O��J�B��������e�`��$n�-�k1��eLq2�{�c��	��~/�e�h�>�zst.�`��b:z��&�v���X�I��2�����6�G�pѢTJ,$�ޒ��
�nD��Gv�ۄ6�v^�U%i�V({������FO?"�w��k��0{F�f*�Gƞў\2r��3�ܱ-I�'J����x��}
3|�ӎ]��8(b�.Ě5���F486� ����*�+�i�n!�-�f��_p��+QUbf����w�#����KYYBMGb��+��=i$6ݕ|d�U��7�:/,�݂���h�>�y~����)�2�.�z�0�Q�g�;	Xm�UZ؜�v��ii$��s�����vQj��'�����툌m���'YZ������\p�`���\࿴6iE�ɯ�P������@�4$j���J�H��*�R�̊ނÛ��K���g8���$m�_�����(ͨ�?�z��@��*a�U��7|&m&���_��3!v����;�Q?Z�鼫�OK-at ��ʅ/ lԆ��Gt���Ҥ�u��y-�`�쩓em@g2`�Wy ��|$g�1����&�v�r?.]�I�Př�Z��0�j�64�C�d�W\�b�}�|���8�@�?a�4x{(��`�����#�"���@U�����v�.�0�Cz<��A��Pv�V/�5�7�Q��r�t���K�o�i�/���PA�O3��+ME��^P]y��	W���4`!��j9Aq�.]��B��g�=���քG�5��C^F�;������U��#ʲ����3�7�}���X��4�F�q�C:o�_^��/��������v�2]� @}�a ��2��YM�ؼ�%I$�cky�}Y�+^���J��O�l�h�y��~�O�V����e�$a��L�����	�6"^�{ZP�M�DY��ٳ�2/%\��hZF�SOa����#2EI����}U����%���7e�3���:K�����zEKY`��� 4L���D�eW9�>qb{Cb2��g��^D��[� ���UZ()�>��"-$�P�Z+r�H���˳��Y��]�u_z��.�Hk�������I�Έts�+���:6:SdR�Y?��V�.?8�z�h�D��E�mH�l�c[�CA+5|/����E5{MhE<H$�LT��t���[��2���a$���>I�m�Ѹ2Ao�A��c�;ok�_��ȳ%IX���7[�i�Ub¼M���� 
�2�TbA��;�����	���-���ht��o;�&��>z���;�a^�V�*���t�ȏ�ub�q��@3�-8ٷ�´L+ ��p>��<�a�?#-��L"Y�N���c��V�����IGȁ;�sp�P�_�nFt���]u��_~� �>��Z�j�[��P|L�¢�D� ���n>�Ȳ���pZ4|I��^�E>�
g�����s��y��z��/F�����3�$.DG�M���.�9�Y��b~����M~3:�cKh��"���Ӡ�,^;,��N��h����Ҧ�ZXSн�~��ы�c����UO� �x������2���b얥�5���$��$�~9���=����NG���C�{�l�S�6�D]�b�=��²٧
t�L�$Y�Qw�.����YtOC\n���:_�)i4DF���zF�n_�0�|%�t{k��!�mR��k	ⷦ\��%V�=)Y.^�V�θ�x�>���ü����T���̓t��n^9��Ϭ�}zE"�l���^��h�^�}�'k]q�}m�x.�^�w<�&ݶ#Ŭ�Bl3�V��V@\Q"L{\M"G0/+���mX��6�3+׉�ɵ�l'����k����a�:�MɈLZ!$�"'Jd��f�e�+_>i�����q[s-�?0�|i��-��9M-֤����,��4R�5j �6���e�������2@�ۿ,��je ���+J�-mG�������^���^�;tN7���AG�'/������N��G�pt�:�C��~��V�r����������Ay2���)�%=ZZ�Q�B���W�RO��=t�����t��6N� �Ib0�"����=����&�)<\L����"7�c�[��c*n������`��_Ro�2�Z%��֞��3�o�9�6��LS3�6��'*�PZ���Z�h?ȅ�;���`���$�.��(Q�i���2dw`�ʞT������T�ɣ�
_ɔZ�t�Hk_�i��>8e��U�4�6w�D)�-��Cl�)��U�Y�,G��ó:p�!���!o�9���_�fz�i/h���p0ǴÍU�c�F�*�䧭�%�'5�OTǛ��G�#��)��[d^���y\Ǟm��L@ߔ����a����6�wW�I��ӕ6�Uhb�G���_Sc��<�����I	�!�.J���O�Xc�,w-(j �rᬓ�D�����=�>s�k�س�J��<R�+�kYi��\2���噮�e�uG�!�"������0��%�a9]��J#m�e2�S�0�4p��C��CZ���u"[����n������!����oH*�����;�����Lz9}��ZE{����{\��7� :�3�Z������%�T�g�x�,q�*ݑw�\*����!�Ћj�����Q̊]?e����@���;V�"�z_��}e������ͦ�����g�fȓ6"��U��H)�{N����sr��Z�<>L*ݩc���]{����٤K��{�.ZjS|{����LLI���M���y���Cb"�cCS�5�k&���uu߇Z��&�RqӍm��0�a{#-��f*�>�YHL�=x5IHl��d�s#��+�^r]qOi�e�5�̛��N�Q�==�x�5��L��t3�>����:��v�x��9��2���M!<�V^�#]�&d�~h��W5 �r���C|	\��1#���ҍzwZ���D������!�`�
�q:i�0'����ހ��&�5��9�L3�{�M�WoZ�(b<�}x��I7�TOM/9� ��9��w���S�V�c����� tͬ�ge`=1�s78�\G���s��c!{����$Ψ@ ��Z��Ue��a���^m�0)8�L���GYq�#�/p�[9��!ქQ���E�Ħ�%��]�]q��$�������W�b�E.�VH�}��C�]"@����'ZO�Z{H�YR�IO�V��TI�eʒ^��mpu��ѦU�t`�\k;����\�Rer�l1�^'���WB,�P��L�\'Q��x�_�k���8$�0o���[�������>�-cK�E��B~�4&S#��L\�r����``�I�ͱ�9�/^���nRk���sf�m<�{�h�5hբ~�;`�=�=*���z�?z�\�F�����?Yj��gj��+����۸+�-�}RS��"Z~U��+
��h6.�\�^��K���h�P�����c9���+��:��㟄�@��h�J��,��e�W\��1���6���r�����əظ���HX���H�T���9hyU놟�&�Pi�[n��A�q7(Pty��GMڅ��^E��w��{����u����9C��6Qr�H9Q ����y�e�a�ɳ;��z�I����\�zS���F�Oj���@�/YScC��I�u�$��e��_ ����'�SrmZAl�-7^�a�����,೨I �����e����l��vmFl_Y�j'����DP�畳�{-V)�-�x���.��.��<ڤ:��7kf����� �5O�z�� {���&����P�zH�H����ۉ�H�`���[��߯�I˵�`4xM���c�z��O<3w��Lm�P�nWfxĲ��k��P�sE9��0Y�J���Xc�fֲO'5����0��� I���9��W����� ��3AH�Y���eLY�Z�?Ieϛ�
��H�	�`�S%�������[
V�����7xt	"�S%۲�W-0١ۗ@XƵfU5�/�����5L={��#�y�8Q�9^4���C1���#���?
5^�	Gg�2��i������/�%����ڥ�8���C*ܰ�Bb��c�e���޻H��=J"����V��IV�8�B��R#��z)�$�l9��,���)ǡf1}���z���������N���J�緪�</�8���t���%9>J�|U�_<'�1пX�K�Q�����{�w^l�j�͑A���
@?����p^9���O���D˅!SM=`��A�+��\�z��qn#�?��e*9ƃs5?��A�le�=F�͕_+.;�K"�M�e��貂:�>kr����={����fP�Q���肌,�- |s���ÑɁ�^�I��z��}��Lc|LL�D8�N�����;X��I%8�ۇ��1�zq��߾%-S|�)�+?��x�����f�Q$6�I�eG�ሖ�.6~�����9���������K�0��SZ��fĸ�f�"#M(lN�1����P����(�{?��9m����|\�(�Oz����W�X���CR+M�qQ�?2�����f�v��{�ۈ�<I^FU�8q!HP�#��W�.�z�c���x��c��[�5RV!�K1� �lP�P$�ƴ5��'��qI�\����� �*�/zDW�Ҷ��M㷊�a-l����H����fZ`	G�'8hK�+gR}2�`r`@~�JuM�ۥ��������p��,�0	�Djk�4L���tù�
#����ֿn1�|�M 
Q|U����Y�������00uˑj=֌r6�a��!eA��W!�gv��V���c�ݔn"�ؠ՚ē���3g����=���^Cا�_	?u<�߮��M�Ѱ��r�����Z<��z�s�p����'I�M��.��e�����$��W��)_5�w%/��W��p+^Ή�Jn����|�o��4�y���Ɂ�� �W�ae��1h�.�ʞmSN��Q�����P�u��1;��tA��QO&j���^zEAd?%�a�IjU��Y� �R�>�.��ѐ$��~�e� FU��ABp��]��񯟀�k���Ω-��R� J���SqU�W~�9(#�E����j���1h�#��r� �%k�m&<=�GڋqYn��3N�׷��sE�ӛ���yo20��'�:U�}���i�o�TMK|-=O�Y����xf(��;-��HZ���W�]��A��$mw/�F�EŢW�%�bsWޙ��W�$��wu��P��]^��y�"D�Д��bɁw��\��=��u%+���ni�i�8�]�T`��1�&I��񠰦���5�*,܉��kA���|��*\-?A�3F���<�m�6IWx��jk"����m��!�Voh=\�R���X-M}�w,�0��pQu�C�Un�P�Y��	~�W{�������d�!�4���|g��v	�P׿֚&�����$�$�|��&!��*��p�P>b�eM6Y�e����;j�������m�WYD s,��������]�[�Ho0!z�6�t�e������`��whU�K�h�>��)��?,�x���V�'Q�CG(���;�rE�i_��3@'}��R2�-ۡcHzi����kz�5��Ϥk��V���ޠ[�SLu"���j�y�<{�>�Be�I��$��'�Q)��C�j7���욦`
Xyi��5Uy�	�5�v�ݨ����ˍ(X�r[��{w+�/ft�O9+��H	�<�P(i�V�hj���7	�������#�����b�|؂W95`y'�)W�U�C`mpd8��s���E� �4�c͊�y7��p\� XS��k˕�QG1,�g:Oec�H{�������x�~)A�V���V�Bw�-4+�$��t0�U �;�,�*|����k�/CC�\�Z�,���S�yb���T��Җ�Twe�6��壩(m��@hcf'7>�L$+<�UB[�dA��d�@a~�0��y�нV�=]�֮]��h�%�����5����f���i>N��z+�4%L�26�X	�|����d9޵��W�`lTp�q�#�% �qr	���`�.�P�Ւђ� 3(@�w��OW�"'D%F�ETu)ߓ�
E�"Uy���k���.O��*���q�		��#��=��V� ��):(s�QƆ��է'gi�����o�*�mZQ�Q^8�)v'��V�%��qĶ�,�b��ʾpjk�c5���Ŏ��O�e�=3u�=�7�R=w�7�ߤl��e&\��X{�i��CPt�<���f��2[�^�,����lY�*� I��qW�3��p���_
����]gP�=_.��&�t3�e.���tΙi���<�U���sL���mP�+F���@�~�V�GBC�#{hk���c���[^��3�6��9-P5Ňz���Z���!��V�^�v�i���qA�w�������l_�b��z=�a|������.��0[|�A�?��٩ݏOv`>L��/�Q��k������.d�/�����8�k�͑ҝ~�_���(4��l����4�z�Tp+�=N0�
�F��$���`��J5?d	t�W����A,AG��+ԕ��ޯ���/�l��z��J֧�.<2��}�����~��]?,Q�1S):{�Ԯ#L�y������9.!J[1��=?0�&Ay����_��2����{�(F���Dm����9%���P��ǌ7�D�*S9��h*���E>�C��u����ꝫ�&���Y���pfT�R�y�2Jj|�f�֛�����K�T�����8̰g�vt~����a��Ȃyq["�r�b�7~[�CrM�*fn�0����[��N�:��*0jv�X*\S]���e��p �gX����bXc��B�J8�wQf鯀B�{Ǌ����< ~4���F�ng�t��	 �N;�v��,����|�͘����^痱����T���-��e�vŚ&��\NE{�VH��$��x�a�X��˞A�e�)�Ӊ�;֥{���O؊����#��C�p}t��a�MlK���yĤ�hL?X��5c�p�h�������?*HĪ�:��a�ń�4��չ�eC���L����5�!k���l��(�s�2)�c鶶 >�ܥ1n�r�g�?]�%�%����/�=9PR�r$o=��1m�����^�̣"v��_W��+�z�3Z3/[�C�j����)�UXa�)c$D�g��>�|��� 1&��|�$�_���o�.x��CYa�]7vOZ���m�<����gn�|�|��X�~&3'HP�j	m2N�f��誌A� ��M�"��\; �P�E+�x"'���ژ NL�����Y �0Q�,-�vK`��9��"-M{T'�<-��ӽ��M�ǰ$�&���R��\�|T�φ�sP���;�T3g�^�P"�vbΚ�N�9��#���m"i�a\��E�8���QcU�|:M�iJ͚��ҕ��ŝf/i��z{.9I���R�z[�xq�4����Ed6[��f>�S1RVd=�ngdI��x	��z?Ѥ�� �Z4�;}��H���|�wE|=)[*O�rHvv\�[�������8�8���eFo���Iw�6�9�J(u�N��uuJ�;�����^ka��2;D�y%|�_;Rn�v���Kp����G�$]�����RGȶ�y3�V�~^�/�D�Q�2�#��/6�3�i��FT F��1�,�AJ�xA�Z�����og���j.ܟ�n��S8�D���H�����ə�<��>_�j�T�=ߜv��|>{�.1��U�����<o�L_���a��c�CN��^��VY��$dߛ�l�,�s@�/쩖q�g��D`/���)�D�牙��ݸ�����k���h"�7R���2q�Q�������"��.#Rm�Pšd��9&Q�p/�rp��~���0J��4�?��3�.�^����ji������0b{�J{͊s��k�����9�_���ڷS�X�)KRv1?,3�Ҋ�'H��nKo��Vʡ�d����+7ɼ�0?�W3���P���r~��$�.���-2��K?�ս�?��b=#5u>(����
���w�*J�:��	k��8]X�W�g� �[gT�'��<�6SY�`��kTtc��A��׷%N4Kt���DV��Y��N�E @���b��jR�H�;+�S��Gz4glĎ�	|E�굍n���pB�Eh!B� ���j��CҹM,�(�7���i� �3Rug <۷+yD�)����+��Z�аk!�������KcuZ(<��&�I���/�nP�� w���}R58@�N�o�x�e����W��F"�x3�;��S��$+��2V�.�yN���`�R[�>(bT��L��6mQ�]6MV�4n�
Jh������u��%ƏLo ����t���� �f
�y��P���E�[s���sElfd�9�v�_$���z�50�0W�<0�TzAR@*8J�_���j|Z�cp����QJ:-�����8�8	�������T��9lb��"�޿r#7��:���w�m���?�WO��Nׂ�4w	J�,Պ�K�:F��&��	���T8� W��wB9�5蜁�l�9� ��NL�mY�+ܻЛ�KcS��{\�H!��j���	y�e��0R���3��l`��]����f��\I
ȵ%����;�"C��L�o�cG= �O�H�0�$P�ۣ�lރv%l�Hv�:��ݴ�
�𗲨o��z�^`�p���L�C��{�Er�w��)��g��q��{!���d�]wpUtD�kd��q�#�{�cۧ'ob׮M�.��?V�ܾ�m�^O���i�ݜ���j�}F�3s0�N�m�K�}�2���Ռn-����;�M��:����!��M�f��ב}��u�����1fLShHѶ���2+�����u��5=�}����o#� '��ֳ��w���ւ�&���!yse9�e����!JrV8m*L�>�ieW��H�Ӓ�ܟ�J'R0�wi��F	��h��@>{��F�(��M�5�IO����S2'�ug��1IY��BȡL�H�I^��qs���A�p��;xH�x�G@YHR*�E���TC�d�(��#L���Iݶ噽\���Lw�� [���C�4\/���_m�=٠8w�J�����M�rӨ��
_��u��Q��Ĳ��?��a|�+{�k)��P��5�H��j���d�>-��-@F%Uv���#?��;�%^K���\��NU��v���K�ciՅ�f��xU��J��b�3�$H����s��0�߹h�~t�)dGc�(��=�!sq=�@�5�5��zڤ���Opf�)\nϊ�a�֚�L�1����>0S�C��<�ہ1��nᦖ �B;]%xE���{n����U��랓��$H����{�TNض{t�����a\�4
D6�"��P3�tSn����E��zD�Mҳ���K!,N��V�������y;|��8��fH��m2[�϶(Ͼ���v&���R�R��@�&qEm��	�ʯ��b�ˑx�|,ϝ~��S�f���]ek���s�O<�E- �����UU��v3�}r52�+L��O���?@�մ����3VT0�ڪ-~��IJC��V�bC�	�L�7�:W>k#��&�0��d����q=	�j��csJt qp�!8��Њ�]д� @�^��q��a T;��$f!�|f�a��`���֪�~�Jì՟�:{(g4&1xXXI�k��y���(#̻�n��JzCE�~�<߽I5��#���Q|�0ͩ�~�<ik�*��W�X�~�h�g���@�����<��gyO,�I��3��x<���Rk��^�C���_����v��)��_;�r� p����Z�{4 S�w�F�u�c����LGz�6��.�O7c��G��;�rڔ��'���N�Ulk�ۋJ�N�%pFT4 i�5[���]���5��m��)����UF�u~WH�ZG鐂G ��^l9�>�(�����D,��k�T���
F!a/��\��5늤�-F�s���t���C
���UX\��W���7E�
�]h�ߘf�1���{���>�p\�ǜ�F���:C;I��T[L�D��Z��e�7g���^F8����N�I�g;�^篞a�b'�g��A*Tr�|ċq-uy+Y�}�[�;�,C��8E^�)3�v:����*2+vi��f� shֆu�*{�Jz��d�I���Bc˙3>Ng�A����ϝS�K^�^�:{G�X`x�`�^6�LO����[M�}u�|�ς��}�	�sy��9���]^��>�-��S��� <�@j�Ҥ_e�+����%y�P�������5t��}[�'�,�՗|�lL���h�p�Q+���y5��!w.���)]!L���bq�i&�y�f�`GB�H$$A<��#���cY���Г�����8� �Ht2��ْ����O'�ɝ�T���j���z��ʹ�ς��O&���6���ǅ^�S.�5W�����,�@��򤿛XNy���X�w��g�H�p9���֌��.8´��/����|����WwRb-��ؘ*�:��E���MR��=���]��38����tPy�y&�,�0�&�����h��U��V/�\TB8Gb�6"�k�h�PUJ�7����bI��N���>���`�t 6dtk�o&�0���J|���t�-��θ5�����!�syF�t+Q�&�3BZgI?Y3DT "� |���P3��Cui� u֙J��M�1��@���f��Iސ�^B����_��N��y((��͝%����4H�ȟ���t���������ۛ�����Z���KB�:.�D`���F͎��̕��������2�>X���=��ۓ\v�,���m���[� ��[b�����I}qǬ���T�9�� ����d�aP�$4��m�X����)�������%�dI/i4�"�O�7'.o`�_O���'_�t���ϖ����,xԨd�$>�b���lf�I����;�P�^Dr5g(�n.���ݚ&�rxZ�=�k������Aa]��qPoj�!�'3:ʟ�����峛��@��.���N��8�t���\<?Wz��881R�{��6���.������ 
�����
��aА�7����m�~��^f�U�q�Y����l�����P�=~�M^y�f��jU<��K�\hƀ�
��?�[��K�'E޴���ȱ_��"U�^�S|���ƪs�w�1T���蜩��_41�=�Ľ�W�v_T�!	���H�K���J���7X�dVR�D$-8���l�v�$~F�)U`��?��Pz]�ϲ�,��kjL*$���- ���	�Г�-h�H	�P�m�������^؉~@e�dC�rk7W��6c��9��ͽ�K�?�
�O��y�$���y WxF3�I~���f�<���ʣ�/���d��:[z��+d�>m4��t�唣8.QYl������t8�+38b���m��1�Z��^��H��n��	����Z�D\�ΚmfjZB����0�������j��$�>^2oB�6,���mu��=Bc,I�����K��A��Lߎښ��S�r�Zm����;1}���f�YeN���v�����;
������A��>��n$��p�-���A���ߺ���$mCϱ!���ە/S�����H���hqX{�^�H��C_v���ہ�+Oh�,wb҆�?'_��v<�\f�n@�H؄���R/�&�S�)� HQO�Xv������U`7�ĕ�So
t����aĩ��.����L����ۥ��&?n�U�˫q��C�ȹ���Ӹ���*�`�LCu��{;�,)�Q�4��+���q�w��_c=(CY����qR�kٯYZ=&���]*i=�����KGN4�O��r�h�[��<.ՌS_���u���B�/�ȝ].��Ks"�����'�i]���T�~eٱ.t�q�Ԫ��<�*�c��5���*}M�R���9ye�T��Y�<���"3s!���I^��8�O����M.��^��I@\*�/J��vꃷj�$�X�3S�X&J�{AS9��z[�n�$,�Do7��w��(�q�v��8ᎄ.����GM++v=B#:Vq��i�@��VeQ-c�"���U��T�� p)憰��]��Ti�/aH�N�΃�6zYf�i�Z��?���zӅo�֛Gķ�j�Id{��2���2�1�~�t�.'F �2�Q��;)�j������7�����&.یB���3���GзL�I�`��8쁪����U�	��*A=�:�=���-��������x	�5��䨒����AmTOF�����uAmĤ}rl�syR� g3����u5����n�����}Gh,�t5���v��¶��@݄F�vW��Ϩ��%���mz���S8�%����MD�f�\|�w	,�����:}�����H�srGR__%��č�4Ɓw�r��T��}�� ƀ۷��3�E��NV{�$,-���7�%7/�wI�	'�����E���(3���l-����H~X#u���A�,|����ךd,��I��a:#^K�
�I�F��� �8�:i% ��շ~O�_؃X�n4�ث�Vyx!�m���V91wӔp^��_�!������z�4�OcC�d�["d0yRP>KV:�V�cLo����}��N�f�4~���JBi��.m�W�E��|�҄{hn��*�cF�L��X۽���h�˕=.��f�}YLk*�����@�H�i9�{��$m��DQ����\ B@� ,n<t�T3��)��	C�� �B��C�tJ���� AOM�~�����:����F��|�V�8��1�h��C�@x��|�F�)�sc��n� 3��l �����\<�O�k>~�IUz�ĳm,:����9�(]�~.���
ZK�Hf	rBYva�&���e�Τ��0�^�9�yG����u\��s���HN�q��d�]�(P�������))��\|�\!�N�0e�Ri��~���ж�w�Y3ŋ�Y*�o:׫���*,��7R0p��mǅa��=����;�D	�9E��"�&t�ZY�|���_�BUou��F�%��d<��{5r_�wz�s�sL��qmЪ���X�s������n9�q]T̪�I��1�X]�](�Gd�.J�0k�$�wݛģ9m&�,�.5��q1X�'��hcߪ�J�=�G���2;gZ[Q��:���-
$%�<ڷZ�7ק����Ղ���W�;�X������R�.>6��o3i˛��ؿ�3��[�V]�Y�gƯ�&�T'��|0��My)�N�Y��&z��9蒱��(�9���XԤ["��vc0p]��&����'�ςd1,�/+�`�|'��0�]ʧԼ��Ӯ���[�KOL�وM���Q�	��E�~���~F�qâ�e��2���0\�A�]�g���~��F��x���؊���
��1#_h��^�4�_wp	Q��� v��Pkݤ[ ��oЪt=-+�/����g� y�E����ia}��0��k��+!��"&�yE��?r�xo�-KWEu	����u�a1�y�bu�S�����3�'JY�Y���a��N�(+(����r?��v~�Z��xQ7I���[@r�ԫ�r�w0���E{���X�.��EӼ�8�������Ԋ6X�k�5N�@&7ZG#�<�z�l�1��:�?T_�9Vt�'��]�~��D*Uf+���J΂��N�S�E�e��LA�T!�AΙ��=�����Gg�H��Cs��7td��X����MW4���I����Bi�je��!��j��<ʺ��ZI�犷��J)�"  d�բ}h, �,P�O���l���� ��*~R�?�O۲˥$���ݱ�&�8�<H���M��2>��ank/�V�6��&}�,����)t`��R9|�;yp}�P�.@��f� 1���lH���kABil�}�dT���ť�*�jͧ%/S�_�S܎�#��H�I�ec�n,-_��'���Ȍ��*�:�h�T; R2��.��I�H��j�Uά��C��7��
����E��0�6�Fd�o
|�����D�VA��^��o�sk�P�=$O��p�#_�J�M��؛��6�蓲�����ö�����kg@ ]�d�>\?W�A�ZG�3�.�?<:�Ц3�P�j縚�q)r�	N�`�>249il�R�\��帲��qꄅ��*(�mo�y�<�,�І��C�)Vl�A��2������$�嬏O�l��!gi����斖A�n�N�	�4w��
4�KV��G��ZNw���	��9�J~���-Ko���ߊ7��=��D3�m�v���z^*n��=V�O<�&x���ǳؚ�5Ѡ�c{�9�U�����+�?�gp78y���0���?��?(��fw��3�{7�Ӫ��Tj�m�X N
�d�F�G�<@�?�*�x̆�T����_h�=��˴1G~�yȜ�!�e��#���O��m���јH-HS�yϔ��]����g�R�u��k�W:��z^���0!j�F{?����*v��b�i�K���zύӘ3�Ŏ�����Afzj�}��Ҵ�A���=^��k�`^�񪍄�md����-U`�*���E�\�t[U���*E�l��'M���������m�1�qQ
���RK6��x�P�M�1�;�B��Kp�6���Ɩ��"촨^�a`H|��(�ZC9̺D"���6�Z����,�z������N;����br#�'����3p)��kv:�[r/���z-���*PQ�2>*�%�'>�Jk�ޟ�V�"&0��iw9A&�y�;;��=M����@�<��
#�@�[l��jsa�w����[������[�9 O��wlɊqI�Z\J�P�6U�hƢG�U)�$����w������
�������t��-Bl���qS�񗹶iN����@p.gY$eLCm\�����)��V'`�kMOO(ː���P���D]���wi�%�tC$�2]���LX��;��R��q��T��V�!g:[>X�WzD������m�z�����m�2���&Ћc�a0��r
�/�'����aS3O��~��k{۟|�٪��w��2+��`�n;i3�^A'��RdK���6'���m?���TOz>�Ҟ7Y��jcG���Ť��I2�څ�!�1_��*,�s����TːR��+=����
l�4��ceN���Q�ƴ����'=��,	�#�B�o�ߣ����,�鵡��ۆ���)L�44g���>E񢖉�Yÿ?��fm$Fr�bC�o����)��1B�3TO>����=��\5�V�>2�Y*j
�%���ٲ�0ȟX�ٳ.&s�|�?+��<K }��GT
�	 ~�71Y�l��]N��H�;����I�P�{B|&wCphn�m891T�
Y�Ӫt��u�M�K�ӵ��(�~-�-�,M �ۯ�� �H�	sm�9� z��I�c���Dm�;5B�e֑I�4,��=K�i��	}Y�����;��o��Z2�0v*�%&V֠G�,e�f�12��ZCHQ��ܤMJ�!2��v?��M���PN�������%�����05O;�1J$���0f�!z����k�@K��7�X�U�-c�#�+��q`h��w3:�H������G�S.)�S2�P*c�- �V����.	�sGRK��[ʽa���H�э�	PsaLP�Z�p�&n{�����)}�Nk����#%X���Ϩ��WR����xԌ���i�'o �d��#�:����eɥ�70?ﯷ���ӫ	H��\�\]D`Ӵ��'�xY�����~^pɘms�a�%�� j�#�`�}u!	/	�(45cEn>z!6���"��3�v>P�Lk���9:��E�'h�)|~�0zb���`[�?L-�Ts$4�oܜ
���5]/�.3͒:��))�-�)� �۫6�0��/�fu*��l]UX����~���Q^��|h	XU,1��XW7�
���H;u[����>R���2%k�x��Yp����NBT�@0�u~�@��rR��x�B�v�5��u�{#�jI;���2Q[H���:3Z�<��fX�MS��㴱dˍ������<���%�Kx����˫\��ϻ<*��B�_������*�����