-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mHLZycKEn5i6EOKcNnky+uYNHClcIG7xt1t023E/ao6WJ0rJe9aZzQYUZhjBYN5YIFdMvMI7S+V4
RyOk3g617lWOfRm8sZAbanWi8oFAbcq59S/J+G9f5YiQrDF84muD4IrH5LwpO5pocjtFihGKoFc+
gG7877MXD/QQcKxsNOLdrEx5lc4quqjy0pARS66GQ8vytFs2SQi1VAp1VGaDM7je1EGGi2mGYYch
XXCxeaTf+G2oD9qL5kp89ogSrgXHZG8PUQ1jnHQXF2bj/+9tBf9EH1rhfTA1y4MUgeKai1EMyHf5
EdREVA4zB935Ow+pRqwaW+zJwI1LshNM7pTsLw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14256)
`protect data_block
Fw2FJTnri4rjqyAJkZe8IBAndK4r9hdA55Gx3D8o3xruNSm2EDYTYwQ77CM3olKf4HGuOh11YGiJ
C7wtvZPvu8z76LLC+mXo94zTG1T1NiEOz+gAo+JV9JxpoxuVqmjzmQMxQetf0n6ASRraWw+8Dp9W
xkjjREPIi01olGe2BKg7J/F+5R/OEGpf9j0932L2rVaeD44t0SiV2KhgDrqw7cMICJuhTBteK5mE
eJFKwjS0JyQM9Mk7xbgZy+z9+HUuzja8M/dBhGTHWm0GWadLdGdRmufHp6V3BVTzQIhgzVZ7BKV1
/D8dRFSMtJmG2ecScstyirB4OodbKGOhP9dEdQTQHXV2T2acey2LgnWpWIvaz/vlTBzdnolIznkK
fptDYiOSdQ5UIj7SFYL5iiLq8Rj+rQLtwP1bsmFD2BAvFuaU4PnR6kO62paHBEyCDvUzYLigvrdO
0iwjhA+VckkQcRx3y2g2wpI0lKJgX6V4WVhn+o5oBL3D43NSuvQ9QUEvzdsADSrskvo2ewXNcz0I
7WgCTwDvWMMAw155E7/k1yp5wo6pcvrxgTfm5jVReKg9AFdUI3NkQUJF1hAWqON8zROF0HPX03ho
YuFzZ4yQOs88AJgIwzImH3bv/Ay8O4L7kgMuWj9kc3ePOWoMGFRo8LiQEVDXeNG+9QTIZWJ3s4T/
wAyKDNp/OjbQbmjV3tUo+WHJ3eVktkmjlH6x+U4y21ZkQOiWMFsj4VwUsubqY1iIRlE/Q+WWa5Ga
enOk/I/WR5AFKbWDyW/NS0l5FjW953iPGEWs7AG4P8Rgi7NyIwnnDMqCrmNYzyBYRrpvfadn9Eu6
RnhU0noFh3WDGUBXD0IUp4FenPU8qSWzVUKaEEObJs4px2xeZRy8JCVUwlTBXwaIVJKZiIlqu71W
JOEpUy+E+PAVOwyZgnNGQT+EMh7DDr/URP4vjbG5csA0BHRx3uSFf6I9vjv2w99qLl4fKIOETeNn
MDU8i/70PpFtCOcCKNs4yuedWiZT6Xf0HRGcECrJjTTySOZ2NCo3vTT4o+zAaIMWCkGNq9AUKEVM
asogZaOmTtHQbiHgiAc8po8uDMWI1Ye4LvoQb8u5/cvStRo8de9/hA3VMgtsKK8VPG9UykG9Oqqe
BGpcCSfXkofzhIO+f3jYCQTxNFj5mNP3goLByHh+n/STs5QLQjI+YZKYJw63LxL3tP9acUUJDtnY
+pZSCucS/T6EZ08vLxQRtmbRIO3ZCzCWIGeHu6aQN1znK1yP22sFMyB8hyp4nH2P41n6Y1T2L/Ma
N3VYi/3FJwFVzSwJmREwsqA6ROscjIq719X08wtuW8GS44sYBjTnc9sqwX0EaXVmoEFcADSox0Jw
Vzo05R5F76K/u/LGu722JrlzKLuqjO8uZUuSVUffCZB6jfZO01ZvCXA6ml7HYnhZskM9q7bSVo01
KCGUCAGK4IMMuDx/JoytzoxdpPSDPzabPjNdOWlEkqYbg7mkPwS7oNc6/JvNxOho6x/hjiULZBKk
fX/Ni0lXQ+gX4m4DXlbnVSTPFIhkLCmmYOrDd6/hmbDZ6CKy18ccSISpVWa4Kkz7BIo8cw2NTAkX
tb1ubkosjPXcf1phnMVlm6GKFWsV4Ajna/n9fMpgqx+PDIsvMzlOgxMneVIRgGAvjwW6a2FO7j06
7FFESawln581yOr1YZ3waZWP4aU6ueusDt4FCKAEyT0P0Y1mLRIsYkNDpRyXt7nCYcWz4/Jp/yA/
QxLSXMFlWQnB+dZhx7p6eUP0VoZlI+8/uwzET6uxufh7ug7p8xJPIWGyEJQD+Trg70zYegBBIThu
TqqUCWgAPOwwjGC+0KmxFa2XtWowUO7PmiTbD98U77EvcWANJ1lV0gfQyr35B7gHYkiz9qxSPW5j
7NST8+YcQDXFVVFxnSCBuQWo6E65u0IIeS+QHdYmFzZOFpTBy4L9BD9lx3x27lEL5XJHdPKFk4pf
8iaeQWG8QYNIQYlxIG0tOT/y9Drqr3gZuHyUgVgHWADxDJI9HyfGLo8zNDMxQvZYpYJ09qV8xMyo
NZK9DoNcVDRtr7mIE1JtScgKeDcHeKzkhaADxCr0eqWYysxJsY3dcNPXHzy5fTxH/l9wrPMfxJnj
ylR7cAiIQ0EVnfjmndETxKOsdB6dxUrbYosM83p74LY/whR152MV6wIypy6Tipy3jm7ZMyvDF6Pc
YdNw+LcPBwGhozUkMnthYBRBoACVBfVQoYRQRsTGCCC2IMyZvhtd77WlySiXAnr1CTmphgadoDAM
ZdUeQPdxEoaQnaUexbVGYO+e7JdrjtNptXXOt4K1F6Eds19q+zloDAQ/ejhx31/BJLEtluK9bgmI
ss24Pme4T3pOb4XSkPsc8QfBF3WgId9PFzdAcQ6s1hUwuSfmMKV1O4GVO6ade+G9jb1ciZQAuha/
IdA/mNum1YDrwW7BJFzNuFkaJy0e2nTtf2FTdeyXLL8iFLA065yhDmVZxiQMq0mk8SOUIQS/wWvi
/lrPPP06sBpHQ83lD6881Uma4OG6leCIg0aPYOXXLygkT4I2o/ga1Wkm2IejyjWsYKYe9sVs6Ozq
xLx/PHUWlZPaFixM8+Q9NytWmMEVGCTwSOp2Wqe78VTzSEGukAng//yu93CIE2m15BRoonvPnie/
AwW7dyb+cz9EHWBDdZUJB+odWX4eIuMRxfxeeBnwpTs1nVZ/TWRwEhjM2++uvVAtC7PffzIdSx5l
bUUMG3uz3rJVpfxUPAmhiIJDvrAdpTR4NO74q3kf/07b/0ZXQ6M3PCsQIORhZ+VmCe4xHphLdWSO
yq+9RYBnDCLweRzbI2yJy0bJNZFPp+C7a2ak8+5S5p7T4RlzU/KoGqSo77ob+GOTBuLB/uszSbJg
A0V3weMTuqOTwgXZakuD6j7wLUje+7yb7hOCi8+IKNP6AyXd5j9rlhazknwRRI8FxbNHZQ3RKo3/
pQYeXce599JGzJbGj7HiNVef23jEhsDWP47Bo3grTHrwXVPPlzopuNZd8NZ5zI/j3/JbdfN3V4Bp
tBm3/IQU5ZrWRUcg9f5Sbj/yYofL3pFj47r8MXviK+4cNMEx2G9EPXP0U/HZVaz3k+UAtmOCKDBk
vEIs56KdsusyTWRPWfW+vHELbPll+kjpvJXU4sSE7qdVn3bnq76Bj9SSVjHqlj4eMTqmupBGRz5u
nLGU333K6AFPMGxz9p/YfGvk8Ih8Pl/n8Xq4qTovVTIbms6U+w4RxuOwfIe5TJlRY65RXA3OeVq5
URv/W7IjuImxxqv9/Kki7FFq1nE8fUNnnrz4dgJgxMF4Rq3q9pklE5odWokNU8C3x8ft9w0l7xOQ
tyLGkAoJqj57casF+QV7GQv7FeE4+duxCoI3UMVNsftNdUEX7FIBIDKPNuXmkxVmoBxPqqpSFIBA
G6m/sdEdShV5n8DINzFPhfomwrCZwxlj14GWUzp4bLabLc70yh8OCC34HAH4jpHXLOnf7GnDgA6x
teFatnug1ynoXrfKCX5TrfXZPewXn6K8N0I0ZmuHvzkJR7tH0iRwibgF7ygwQOo9RceuwPoerkDV
uaGQapEXJFhKH0xrk2SMapyrLMVvrEXxS5+3LPDouMiBE28wCYfUZ7mim7DHAAjxBfq9yzCJkLr+
z1UC+azgGjXuT/2LwDQ3YBtjiuhRS48zMazx7GSNIANUMc2cUFzX30Ocni9nRiaFPjQVkG9jDOZo
t9QzdXJTILaVhjRYe25g83SrtIV+RbguOK2sDpMN6s0/BwGI76xP1n1Mrvt0P62etviGkQxg0oi4
oKY2XF5Q/YoQ0EVKnpJ2WLnVz/ocQRROZSD8CdoKbG7yUc/1UfteMusxePD8R4N4clxjZYvIa8do
GLNdGgqBH1H0q9HGGXvKXTo2kq1I+lYQZV9UP8byiyYvfivkuuYmlothtVwiyQIrqkci/ZX9ZCSo
yCVYJPaF54NNS7NA+LCxp5emE7CwT+695Nro41ih5bDCiwqEaspDZ7aRcuGlraYEeET/Yxt+OgiN
rHDjHwB/g8ITuERT+3rX2S+WB+yH3QE7cGeW8InL59Hn1nPfYafAkxbltcKRqgiDMTC5AAIDmlYF
J/Xzdk0WrwTJAeV86fm2VKfvCBOr/WiSsaIrfPkysNhlYlRQ0Sbkd05EnwU6c1wqwY3xX369IxYM
70vY/jSTiHoucEQJcrVYWdFCIRcF7a4xPKyVlNnjVvpJnDvBhPpgBZrtjiWLkw3vLh5X3uZ6bMHS
UZXff4ekqmJP55pABAgsOfKujmC2c+sIxpoYPUO2v3ksftby6KdcNF7HFyG5XJpLfb88El0LzzV9
gx8xyXMBmdddSUqKUb8wHwHU4jNFwiAPGhc5qROZDfbOezO+sRe1RpjLdZngxxsWwxKbd/qSdX+d
TjrC7ViDMdD69QGB8X6BKVLso/aOGpMU17VMzq8GHznUTmIGp6g971r80zpMl9HvmCvzOmfvGDTV
xK5vuqc6x9Lhgzn47UsQ5fdyLRZyTE4+WhmnptfgZPGK5XzEEAtNzDFfvsNfKOZidqzuEi5YsPEK
yXBwYGSfrDA986iq457571XcrFlJk2EEm1c6oV/KAmrzKpSWCrukFJXsgNdT3rs7HBsCQh4Ef3Ss
tpZ+Y9D8JH0NvSFxSpifkOYkmGBms2UnbqA9KGDNZdnIEv3fz4LxNA7w/jt5+m0UFvDhCSH+Vd3g
gScnYJuP3XCO+wXR1wiVkISF8QyRDcPf9zbc1gXbAHPYGPMqgc+jQ1whCecqasfLS00TEKQnCfpU
4txPdq5BMJgc/+ssfDrh/QAz8Ft1EE4gNeIq2mTvw59vTon2Uhcxc04XuXleVF6W4iEeMLlA4a3J
a5MH62AhzPffJgnOCXpDrpgqB7IIAcT6+0nyOvyj3zgdFrH1NHuQRXYrUtcHZscXP5igYGrskwB6
hY05I5Efi2KskxSASXIbyrLPRLqlzw0McrS3TxchHzSZUMfdr4N0kmXX5RMGyCD4IIXOIuiUtm+f
EeDGs3RkxDO34lNvW5Q4oZUTXCCeY/jR1mEZ/uA6hzTm9cNYc4LJH7DUnFvUuyuvUkbkERCeTizR
ihZbi1yRDq/HT/nJS+TLugnyMxM87tSy9WIijfm0sLqFkBr7FU7XGOppRRIUWb899YtGsSqRY0gA
WnlmoR1t0/Ln781DoJzpuYVVN5x6K2f//Qojc0TPcr3huuMSNZVuW+LoVp7k0eRYIgtbzH+BGDMf
jCCAPEczKRrdTNpUVGJu4y7weO1ZIqDYTm8EgHm1g7fxUyqnvE8W1nYTqpwKErhLEFG/WC7+DWLL
ysAq//O5mZAoJxbM8RkTH6D1OpFd+PxR0Wmc9UtzopDEKPLeabR+2ErvVxKGmVX8F07xPN+d5HxP
PoPabzGm0RelQnsSJOirTKqTRFomqzJINKg4VC5bB/vqq86dDmUnybRiB2fqGbZcrGezLpbZVtqB
hPUSBgjvVBgGZMflxKinB+Cg82eAT0hRy2bCvUjtkWQ53jPv/xP7ySie5DEfYAyBvNo/mwrpp0Zs
L/PLqW7hPkTG1qA2rFaXdkUdUAjex4fjzl0eHCn8cWix908L8KnjNp88vp/nOnpq3EPeg12iWLJ4
u3/Ru0wYvz4zvZkqHf+AQA8LV1MsiQs66Kw1vef3SnksRbt3YQ0Z8YoSZ6Y8dQMRXo4jISDI0ue1
7h+DWmWr2LvcMefY8iDCrpvsjkQRYOjO3viZ0eafR+HeBjuZodxVn+5gntDD7eytWhWMuvOnPuXL
jimIRjHkv97Ts6BbtusZ5Odah20AeQV/xl7fFK5kxDe7x4fyGoWaGuZ7yNfeMp0pDusLaa0yRVWF
TefofEPMhgntxygLtjxIl+QU+vbnluakOk3POELjI9cErJHBDWfCS9By5UdjZTv0306w8WmJukzt
I3c7px46pfATpcX31NHSF7gG1GVydB/ltLQnBQOjpaFIUYuJZiuFNHe7S7CnbFeq7zMzOU0bAHGr
/CVKoT4ljKhzLl0bVGVp+9bxLris6Fl+DRuxek232VVnS08rEQvL8CzlKFyKNsdx2VTvlec+55OF
0R2BkZOc5+78KQSiI2lAbW6lkOfjWGFujZdyuZGJCiJ2aqaLdrfV6C9ioAjDFP0cMGscnn2P0XjC
qrXD4uLph6t9sgvK9+PzIIXOgpmjgoE61Dj4LRGFcKxumuyy7KgUY5gEBsdMbAPDgxoK2e449QHf
h1xNap1K4inVPozIo3i51SNZHCrkvHdloQIwzgfXMpMMGbNXz+Vs1+dc6p9BuOwrairJA2ALRRwW
1oXyDMBjXVQ/enZNc+WsF3n8LyZCiQO2E1QslLFQ8LwvAjQiCz8fYbAeUIwvTjSPRP5eWpgxfPCi
pEDsMLnO9FIEt1w40nr0YZHDTHgWfHGbpKUjot2EMpJB/+/FP2UMODrkHNV4ZULSrrdip/nGMkxv
O5tHGd6mdFcgYaIK+Ownovpkk0DbsRd5cUhoLMaIslnIAKAhogCOLzeRAANOYu9IJ+i5Y4wpLGrm
FlEM9qaFyzfTQRuGqzZUT2cdip30+3qrr5D0Ec9nBTEX/k9m/qFqPYGCDgOHXSqfEhEqxf3YLyka
9jJUW8V7ORROtc8hLte2PNUvKblL5xfm5W2St8XuWV8KooJ+5UZW7taj2vZZqdqkWfqxmn4HmpOD
T4mVeoBjxT6iy9d1vS9M3732I/Gku+jMRhhEbE+n8w62yQeH/Mlbt5cqjNK3gTox6yVeSAIMxlPL
QQu6n5TKFULwU2Yc8MxDGW3+tlx0kFBjCIb+SfZ6pCIEe+VGioPTRNhFLq7IHIET7tcUeHhY6zlJ
uTwtElMvQZ3D2Bm3qZ5dmfTi4ya8DCh4YkELEgir0TatIkJhdAgJXW+/ePFeTPNvnVK+fjNeF4jP
SUCiLlQmxYtrqVgAkHMUcErVzUIhEsMzaRQgFHZxdkuKRTaBdPD0RGwRruHSKUqq9+PkAz0PE9e2
LOW5ATuWLgezqKU3Cvagb/1A/8poGq23xzfV5kjpr8iDON++XBZS7fDblPZYkd7+B6lSi0AinC82
0WaJjA4lT8FgcZSRq5KXBNyRaRECTW1JuZeJUQWt5meWdi9qsjGSj1F7CfwTf+AbqBZIL9RhWhQO
Kf0RJ30GEbNoph7L3/lzWzZwUsS9eKtELVNVUXR9HQXTrm5jRqZ8jpZvQ3z1hZjZ2RXh40gVzQwO
+EBzVJVtiWBG2o63xWvjlubvupi0RJ+m7OlNgn/ku5Vkl/3UDajjaGTJfbX0U4vQSpZQAojRU/eJ
CBQqNLoECDbe05sR5l0Wd2m2vXaDwRUGtC7FhIHDjD7sRQh27JMahde+gwYFVTGDob+uUiAALJer
46mWKlI1ZB9N4pSPoIIcHuFrQaMJ3dAR0eKK+C6o2LbL0NC0KFeq54K9wPPf/fFaPo9VeemTEXd0
f1eW5cZHBSu0eo+4rxoGIA9YF9mIko3LAbiKjubXXDvPqp3RUMx4ORlkaA7tf+LKyrjYmNtv3AOH
Png5l8ydpVl55WYpZljpZ2auTn52lHSmnzpFtwdHAaATPe0jqwecOqVl5NsHDFhcE8rjWaAVQvZ0
2OT34J6aUcNw9In6jkBkAowIS6QV795Un0tcFECbvqmHBteEsWdqun/wN3cbymQoxL5Z0N+wlPbt
z9oMSfngnIx5u+XTMWTO7K8norIk46Z5PmaIQkoix45IYLB3/AYG7tRbhr/lBfXoRDlM+NuAdrtZ
WYQQQSHBfWXkYC/cIAvfz4bi6zwLGoaarIU4SX8IFUZqYKPtoUsSa8l88cNzGrfFhyghk5wdDdkS
DnBVePbpMBYvsLIjYIZg103Yjfjv5fZzb68A7vYeXULiOkF1+RqOfWwTE9uGp4o3dPhl2vpxD3RZ
skzoATd8AhIQ9M4In1yGO6Th2bG6Rb0ZAH2wrwPoo2YQUdRvkTgJx2V0vTCmBrK05WPYReeq0w/c
mNcF0r/iKGGroR4A63gMO2qNHCSwr3ybODDxbbRZVVa+kEEEK+MOTMVdIr7dZqVxPxQSL2p8LkQx
cZ99DGcwLf+xOZ8xd+p92fH/c1oiiM3ePREXtyAPHWpZNUbtsBJkdrTrwdbhHlarfVxOkn3XipXs
K0FV9tC5A9YoX1HsPmO6sdifSyxURWzeqeCURpXODq2slK8OvvzMGHJ2TxoyyR1lHclI5bul4gjY
HYXDF04WHl+LLBOWLBEnysU27gpLu05VIDiOp5Z5WUqvP2bVDWR+mC+BQwsnqcHcdWF4Pm9aecIa
uPOLdvhIF88PI82RQMytlNPl46ErF6FwogS7P7Rgonw8YPFYp8cYMovH5BKepj4Of4TMNSYVAyFt
rl3WovNnBcyGVvlbN656aEhhPof/hN9Q/fkTYskOAhmcsvKdEK7qEYQrd1zwyeehYvf5L86qopgk
/wRJnCnVzNxrLefFPLgL4YDY3HrTHI/nCNbF//iDQPoVmi8tcIWgtCfPcP6rPvgiY/fcvTM2Gwzi
GhJOzRCmGlEXg95HsY5QijZPniekGLeMPsnO7pUSdW6+aL/l/tqMxL8CGWKJoQTYDwYDKHU0W1dE
7oPWLRqZbSx0nqV09VdpIWFE5tqoMWTClLC23RTePRBc1exWK+gIpaPS/vC59yyDyRIf8Oi/GmXy
RVGMn8WL4s+yzUsvRge6Rs/FL1W7j+Z4jWgDGrBORNjPQbBkqeiGbJLdqaoVzRuvm71FzM59S/wY
+Br7KEFB+gTNyX9pmaHQ6CsZH2Mw6q8qT83Fzrca+1ntZN53VMSyHU8PKP5sxYvXCuI7Wq4qR5tr
dMK/3VDsu7m/VBLPATE0LiccCbqEhe7AVbl7OFc1Z5QL8oj/JC83a3M9tYfuOkpaBqNwMsN3Ai3Q
cvzH3bC+Zzd5vnBUOp76GQz+1K7Q+XKVWb8FQFYNXnjw6JKt+jS4DOREhPlaSKbVkdQ3cwt/8THG
2mPFKlgf5fnsKwcTaq3xPLACx7ao7DLTXQ2D1+X/63O55JnsbwyRo5LUqSp6+OC/R1CFnD8HBusq
2FKQ+4ps3UTZDd7pECLFmejfTgHsqApXAi1V/Vhzj8DL4/KzaM0b2NdKw9UjGFcYW6i4/r1XxKlv
eWoTZ15F4GMoPO/BUSW0WgBJEBOSiewJ6wmxGUiEiH/th0W6qGMhvv//I26o6y/GnJ0WUOnQlmFd
HIwrsBF+cCTVDm5NxQoTqjjVJW47dABjgcjer1kAq7An9BYwK538M/AUBy73JZL21YVIjnmSQzpb
1lDT/zXiDxzoL6+JgivrXpapg9RLqoOB22mS0lO55p1Mg7dAZNrJP25Dxytl+VxdVP16Cp26KM/y
uRYHtvbs6IE4fH9GYMSBaUkyaz83FAsM+bxOqgD0CN5DMy1zMI7NExh6XDlfIo7MKtUBUmZ1kRRN
0fvEKMVyojBCLBfvh1kcXU4AYORM9m4ZDy0lxzoiPl1cdV+CL41gBMzdssg+usjPEpdFk1c7+C+w
L9ULsQyfdNEy6yjBKFNlRu8oFvriv1YbDnwtwh9VhYnuw5AMpQf3NR+XEkzasJTYCTE4heFig7t3
tJNtrbpN+Eej+HRUPCtxORs6yTl3R94wGZBUhU+z/IyYSFqpRnCkU1lzX1CapqioxZjqqKIfU3BB
+PysflAZxDItt6romGC/hc3DLtuPP/3dx8OGxUL9ESJFdH+3Kk51vC1k1uwd827kv0lx39bS1f0O
bjeg4fbhh3m+lAX1jYkJFaeqJRnCyqG8u4qrwgtKwEQ81Y6Zi6fxwDIfzw80b4/Y9JV6UaBGDWQY
qN+T82apQnGNtlKdsPWz5mDRw9I08Q4W+YG/XpPf8e57hxdKIxnBWjV51AQcBp27t/XnmCxbv3bT
Th+1V6wxn7a/tQAoqoeg44Y4VEuf7tMYMFiUVQT67fQt1RjzjHneKUeBQHrCNAD+htvtN2BQkF4b
OXoJ/tqf3lmaiV7R6iY+SS/tzuXXOM0cYCCYnv7Y4o5xbx1qjiWIv/aXRUQmaoX3V/M6ow8m4X28
kcvVECaNGbnLjeHc0rtHORPvhI0BSPQmdMNeWepHw3+5ILOfnoW5s2xofZjTNN1Xix5L1S5ck12A
ar2NO4x/PnC4rmxpCf7Yao7gI9KI5ahvsLHG9doyCiAOEDnS351GgiR9uWN39FAtt3SBtko0hpY1
BX1TiiRXyYZS8btri7oX1h/O8Gi9rMt3XVhGJOmJt548MGR0e86Cy7joHDfWNjB2aU7beaPMh7jV
lhpNywEZlWhVONWACGmexxGlHljJk4IE9S6Sz/YZQvKTOcBK0SESw/koVUg8l/bhnapCVlPvkMPm
GVPqwBhPf78RXzdUTEnrIjdGyraubOtXCgnnPnzvB8PKAhwPNf6BKDhTrdbQABGcaPp36YABSVBn
ijDxp8Eu2ZOlZ2zDKYkPFRg6Jjv/tFyq1JuXOJ5U4wGlWqFyshJJ80uGUHG9arDoz8SLJrpEp/V5
yCwbujTDsZKaA73nWAI6XLlVK23Ibkn3CFb2oSdHMkYGBxmjC5coN0wlXCybG3opa6gkzW7x3ORP
9JR8KAbK0BRTFOOYoOxhrIF/4m23TzLvuGHoMEY3jAQ88RE3tBQPilADFZ0690yy2cZYsG8GJcNe
oC/db37GH3UH63LuJrQf7WY6Mb4wILRFuLelViEtnbAVRN1Hm7Yf2rkQSaNq7QwilG+EMF8p0YGf
leIBdXxJFpkPRH1efLgNTd6KSoNmTHIcnHliK9cbxAOsg2R6MDZtvZ5widM+o5tmSginxa2AKPAo
J3FPo3HljwYoJtVHt47JNxxqMSoqRI8lPnw9esOf6F7k356BJyOi593DHkajzKsPOuw4UarVRD3+
FVFuAgwSQGPAAueb+/zjjjzAf0hAG/mfn1Un6PErc+tOfJRZBZJuORLHrPZIHuqBTBIR+EEAVlBQ
a9AkNwCFK5mQyW39ZYMPOTKkdM5qW0v4XMZwFDT8x8I6gIO0LhMwau+JuyKyMBplzduN+NRHXYzV
k3RjrDsbowJGhJ+X0E1ZuJYkAVPgLKDEuvnQiwFT9wt1yqTH9Ilo9DBIzQGyDCmDWLeK1j5WpW1c
mjG6DNRKYrxZXbkw7x/hxqNwYCum0zusc44iJAwKYEp1vjDzByKzfaQRubm5TBfd/zM18MyjOePL
RXl3mNis4whSp1kU34oH6NvvWquhmIyL9wlWB+WKyIGBsbeVzJeSMUuxkcEple10UW0vMwKrX1/U
AdOC79vdSZ4RkKQSlNMVPTHkv1W+/0p34dr6Oj7R1zXpvH3j77642+AGU6yuFM+cbJr0w4Clq5c1
fAbrTGduDYV86Ach+7yBxYWKIOua2eEmJPzTjapdCuV3CHMpDCDIqVNAa2Mg5W6HBQeAp7CpeWwa
3gFGU7Jve9GtidRGtZQPD50VuFggmqgXZlFe9T8uawe5nn6tskmErDVB0HVuMkFmL7fmILE5rRUW
tQE2ix4UC6mwZtVyZg3PC6pKM3GwPatdfpliDTEPPfWGsSUg9cQwYTfrPfDf7LP+qesLXFmk5HLI
7130jgn4sfPcWbZ+dJIpm/SnwRAwjsTHOkbiRLgLKStZYDB1e6Vv+BMjlg7LmSkzpJ0iu/Ic+1vl
mvvZeJcW7iSKasQtXHwiUuG+gvOKtzdo64PXsd5hBNXyz4GpGtDgkRhR9rsRmDvpE6HYQ4cb/OYP
KnUp20OVyi9VnKzKdtiPUKgADDOozsy687mJ6v2RnqJBsvDJw6ZyE8p0USpLS3YCTSo35Rr2/wng
QWIxM5H+mYVEI9byK3zrnckjxT/QYB3xgZVTQLojqQStrpE9G2NUBdhFNS+EvmZNyYzsIxmU+hJL
gA1nqETs84aysvjN12zYpKHhTZ94BOtYpWgBDyJmsKlrsuvikG2lQoO22U3ulVu7aCK/Czlro9ki
8PJNpjAZU/7jOwBjlJuRNezjKgdnjI1qOQfAktR0t1r/q4JU8Au4EQX7knOBCGpuw2XN1x6iFMYj
xS4/x24tPjbmoTBHt6BETe0ADrNxS0C5XfIIsI3W8chGBwirfgwTdQs1iRVDecs1M/VrRHM9tMCK
hLXvfrd7TCJNY6e1xx6NkhWzPcRmrH1H04SGM9NTa6m0OoHX0yCnaBNgzNBV/K1gU8n+8HIrINld
NGym1gBb0PsMEZhPGpnRFQ1ZuTw2hK8OhcULjO4/xNphnpDez/w+55iboJ/5nTf4xzI9y7WJlQSP
4PpFvdHnjA/5fQSU+w+B+DpjyqtL/3B5K3fb8ElSqU7zFJfPTmqUJSTWjrgvVxD7hP+okKDlCwYK
4xJAOYBn2bS4aDIYkyCM7vcTEyVobjSgpnOFRAprB4+bB3pZrRAhmHAnMIZsXTHtxNgZU0M74yUn
xpV2mBLqOWue8vV2IHF2kvFo/BdY2U8uDUWxOxeKIv70NnliMmvvAkt1zHMpFc9N1JLBjMZpiGLL
dAv3GfLr4Vt5U/CBo8yToQWG1NVlQZM/+i9Xcftnifa7nd/aWHl/bvOh11I3pQSFaEA8+0xtP1Vx
zOfOtUFAFFNg/iWgEV9jY3R0KBo3oL+yDJGyipJWKV2E9jqgT7DSb9QE97JEXIRrxJkNjaJW3SWK
qKwQPukPBv1SAcTSP7M1XxRQF8Yfrx32uxt3bbMHT2+h30RrEXSaUwy/+FF2OpJs4j57TanhjgMs
eJM6qh6VCB2+pFg5D/y/XAymUWYN31t96iF5YV9pAQbvbNh0uYTme60h7a3aG1G4oI77RO6/TkK0
ez9jTK4tBm4Ly5rvCScFqwcNxVT0h8G30IiW+jeP6UGtuLr5NFuJFEkki7TAnW4sg4lH5VvF2r5d
g7Ks0zfvsFAHrRouSNM9uEimkkYmAsQaOgTyo02AKRVLpDL/bA0IuMtfbW5xyhKNzBuqbZ8nRC0e
FfHyadq6Nc04HjTlOQ1rlxoBqdK8bJTZKQZbYhB7rmtxzSlX6zdo9uu1d/cLh3H7NYPFPZH0exUp
do4Kb61t9NQOear/moPiW8yd7nlrVPJi6BJ+nfdqbCw0dmbcHD/OyjDlBsjMSpLhzVaKQ8uMf3/R
+DJfL1+pJZ14NYqzsza/8tGj3Khi6JEv2+sSZd6g+kJ1hJUxIGLaOn1MdRsvQTzRIQ1e/ApI6Xrv
X3PdMTw2uIAJ5ILT6dqq1geTY3KBrha0syNw7mv9mRg+j+3k7exMIDpubfda3MhOesG2/Tfe6kmG
i+/KhSbYxRjzb3tOwd6emeVXUHE7QClqHlVwSgSe3eiEIERd0k2M3hUWH87XN23Z6zwz2HwspsLS
zQROr61zoLEDUHRlaz24zGQE4Ywy6gAazJRarklLMircGtueJAQmYRNh/bZt4GAGWpZyEVlw/2cA
02wDlp/d3ssx3raaCaiSWE8C+AwfSm+KvJht7OCEA1iX8Ln63Dz76T47uwcXGbcyeQrEiu8Kr75J
YQ2ka0kvmALNYcSkuoHSJEJJL7yblxwDPBAuOrEBVPwQbYQnu70MiTcbc5fgFsPJ1iyc06RSlnh4
xFHEMyUtAa2puY4Q0Na3+iJrglfnEbBWiyIXW4A3DN4NlxZF172hAcVV/wD0ER+j6ngDXA6oUOZx
aWE+/bI/0sEXvOk5u8FFBAwDkb0YKBitrBYVNXuys3XHodYZgJxiHOwpYrYrujXNCj4PESJIfX/g
gpZYSbO0jzNus9RGAwJaarn9BlZCImdV4gRXomp3URrU4W2WcLKqW3tma+DxlDZ9Yajsm0IKDICe
bUNox4Qusvc2YTp2T50ZY0KQvZ0uCclWI2bHNWEC7DJUibTfw6rkbv+HQIT7NR2u400hmxlhjXwO
3+pGjIRM0ejaIOiwTp6QPsQXB9FdXW/0ZSJ4voCPLzqUpZ5ERQhdn7kFpuO8tDokIqA/3BCqZExo
09ejAMwXYGDSEtI24pcv8pPOfuBmzJUJpdxBdxjNgjSbLhfsTKYmNQaablRKPdyJa8FKn+8bJ8lJ
pNtgNy0yfd0SS+rdLVR2BUAnYIyEcycBGCCZkGu1b278+bjuhAF/wCrGsirfEmSxbstTujwHDHXC
kaa/3pkZewGykukir3I3o+29v5fXk4HIzj13vSDYsOcB0WCsadUN8A38iQ31DrOI2xCJT543JlzL
wfErex5fK03SbO3QjVW39V7v6ijTyEvFW7rUmuqPIApcmgwheyyWaDlEZomvY4F+bQtqTce4NFCu
wqLd1JuonBn3x5JMWvtez7qE/5ds3N47RokpM0XktIRGE4jyUHLg7Qg9MjmLsJC3wgH4UvqPm/WS
LwXvYHqN5GBYsiJhqj+1EqQlCQQzbKO9A2OWh24Xg6M2LcyhMwcnEFetR9k+E5Evmszj1NCRPpbO
tcB3DyLAJGi2VxNuj9C67GZz8foBjLFly4iAZ4rrqgnZkeZSrOGh8zAcastn1rafCMitx/E/JLSc
McifBXrtcOl9PutDHVqp2ieF8L4brV9RtO2Qcr4hdU6vHjEZmXE64Cez7/iaY2nM5aFgEL3vQlBu
hZ+cN770sR3K04Y3Ujpj1Z3K5t2k3fC95GGFZzK0TISctL2kpWmvBOzJHOMCdoHGWwmrY9hDjXfT
j3zFoJXgNtaCNqM9LZJyf0g/KcshbaZdwuBb1sUFUyNe5CqHYSgTaedCDj6YSdV3JhlSM0rQmHZR
Wjsf0ARwjjMcDvPtD/Li4YBkPvHB57bjIhfGOQ19GR5o/57YqE9gVkb89LbFOHLLBaOqITz2Xt0V
eqKeoDSJTDubvYEmdmi43ds5Of3uZPJnrou41rYxLA5gizkPKNKzyTdMd3NRlx4ok671e/7oBgtX
Vn6mDAyHHnW1ndOUUpryHehJ74ivuVhirL5y1ZDdosVlhbirupR2VeiIo/Oipf68lnVr7/273NI6
CxCB8IuQuMKObyDiQ0gWja9UvPYn3RW6wh1i9SfXLeHJ58xeE8yTLpJNYNREnrqxJpNogwr2RmTQ
YxaCe/P+dhga9SoS96XvmXQsh16tSYur2+bl+00Rrx6Eg74YDm4ieagrJLA2ZQvJu3NhkkllVanG
4QWKUOUXsezm89ofPegi+4lhKQl7EIWsWlwYQGg7TmMv1s+VYXPVF+/ihg896ACrNp5m7iPNAehS
NNyPKfhvC6q5cKMMPwStl5oEOm18rJH46sRxJlOSIZ0yrv8n9qIsfVqN0/2cltPN2LwlNVUVK0H6
iEm+uCdITYtzA+J7VVYBHyKYxY+iom1sRryhixoc+wkgZeYRD8ufUTsSOBavHwe+qvNj9ONq54Ie
iqJLdrb5QHz3x+n4uiGQgYDSfn1A85wqrctezFF2yCxfvyUujDL/Uh5E1ZA4KnZZqCv9NcNmlmoy
gNx1UQ2rbcOvtIWOWMPAB+kjVtNJPOa5k/EcISEqG/AtibtonidXXIHWI3Bd/hfrZ6C5kdpXI4B9
CvyTaI1SqSgDbO3DpsD9uYSk7Ack/lFspWPIgQ/Y/L7cTbaIq9NhRIYneFiK1ZYIvj2biNKbg2Nv
HwQzX4PBj2QLNtlrBQ9/QjC4k6buuRzbe68GETHpkXUlk51y/NEZlkgHeADxWCgY8gMDVKD8srLl
LI8jiCYeP6ZNtL+CJRZK3oZVGJ7oglt6+KTxVDLatb9IQ6S01XFoLWbfyBzCiLSGbLMdqLikROz9
00FQvFwDjY07Ts19AcByfMMpUHM9EdDchTk9ZMnYJvV+nOp2UrLAg/85xqHm97wmDzvrNhl367Sg
KpYjzOZp7SbwklgDepfNq4v9de9VJpsJynHmRyq/Wjx6WmGe/ojdshOCqQ6z6TM6mfukBmLYrvdn
cLfv+1Qybbpfnjp19lPHogjsj4vj02vPX3YdmfgAllxa/vdIoNCMw0WsgVFMecfrAu7l+u8pIcJK
j0BszQuOvAKoLqhF4LsembhhTYLkpl0M6KP6nOdc1Lc1wfLUna8Yo289X61Y9fwzVvrI8piAiExk
JMZ+S6nxy7Afky0E9ml2ZXq6MptgGfps8rH2+Hs2KcCXjBD+rB3vNxOZnYuRRY/GqwYPyYX2mr6u
64FXlOXTutrfZ0Jh/4fvOLmFnk3Or9mcqWZzEyCyEEZbE8jpTyLnWYQScFGo0LyB6hbwZHOXOfxa
IA7ORaZjQcFl2CoyjJvkR7LBQ1naOIlg9XveAA82sam20YLsBbAzfwH2OT+QCUJafi/ik+2i33Ui
+pg+uY4h5VAoUWrg8A8ZmSD4xeB0No9AgegktYb+XpJ9tgAthIddnQKDhLHpnjgtlr8gMJTLgUtU
+HtLSmi3GXwK5gZF6aqVmjZqN3k8fUGA46JeNnB3GU06xObVHE174ImXg5NLoTcEFApBFz0omVDw
ZQNdk2Rs9ZIe2SYCNAVs2Pl6d2twSLOMOZ7aCrrLgUUAxYi3hKWAHIUvQhpcVaf8UEc/LOvJk0MG
C/bFBFRudPcBKbEb1eY3rBAuSSW4PmBH8WT1HBBP7smM/LkqJqvz6W2OcQPAFYRAu+dkw9GbPv7/
ZIhXmQzILHUO6tZq5fjEShexjIKuvVRK8UovedhQiWxPMcTrBJ130IiTGS1slx+B6SS1kEVB9vqk
C6qnpq21QvQ4kXuzo5nG4FvludIgprRHrxDKE0d/ZpLedIx8U/hxL2MNN472SVfSaq7hXO5oEYDN
u2Kj0T6B3M46QHSBf19yvdpcSPnxQdDdMz2YOUKxvSXWFTwKtzCkcN+C5NCn3X0NX/Pax+QmIbUC
xrBY0PnpBumSeK3dxyEwa7CC55TxYDV0Z89Adj/32PngnQPtiCNWIRqc2/uq/nazJUaed50DYelJ
yrmLgtuIa0U+7N0RFf68sL35RG5WmFL6Ve2LywRl97aXXEGEtvhfRgMNaIckvgWk61s3BQYfnVcl
4q6DULiicpsfprM2SdBPLfGWNWv7mX3xeYebuSnzQAIxqrqa2Z8IdDaSSLisoH6ueGu5POSSPS16
NmiW8hpQigsQwDFl3qNcDMY1/uLc7JyWPMwUpy60U0+J95Bo5f8gPAPPDp7oEBveQTNDWfBk4TdK
pDA6UVVesOOlN/UYESrkgerwGFryKFhi6B0jjF/BaMy/7eVVu/Mmeo1M6XwZxbbQGt99yI+ovsZj
+udRhwgmZ5Pawi8mhK9vpw2XZPmY4GAIjFllhVFBMHV+lFNJEB+vx9iKK7w0+W/x9rGaICqVEGVU
Mw/DpO6bZ5Ri1F78yAD1Af9IXyiIxsJl/v/7oz/nf8WXgfdihO31dzKFBJKpinh674i7r245HOFK
MPduEImQD5/xHsYhEqJQrkvDZajTRijigLqQdnpbD/T8I5aRYBXyC91KS6E6LeRPUkfgWctHpvOs
6JBQm+/emt4Q/8GdotZihx3wYo+Y9wjQw2+cBQcGQiAHRj2ck8v/0Rt6njLhp/BJ/RIYwPLoKk3v
4wsdx4OUAKZwK3De1UJFqrKl7a3VoMNZ3VvWRDjkypbyJHVqOxHawewU+IU1MCBvRqT4RBEIj2ff
f/stRHIf65q5FLcPaHj93peVveXWvl9Vl6bSQZ7v1q/BB5BSzelXEm3l+/eoAMY4C9gAaIXvVrxv
RpZSw2e7I7BqmRI5egxhJzRATelhKxlFg7fIipWw9GFFS0YfWoFgQc8E43fywa9FglZEKiSLqAYp
vW4daL1KMH+F5vRDQaWh9klaExJwF5SKvIcFqGZzMaFFS72Sq7snVPN6lU3ejXpMbBvxmXV5STbI
ksMolWzJyGx3Mxvi+hui8WSQTZjsQ4Au2WStBMT3j4IXcngrP/ilnAVVr1LLrszs5zJszEGeHVRB
l3TlNkTm4iElVpWVIeqEbR2CQh4mryh17BK45o9Lm4EMHpe+34JJassxTSFVHgEfj049GtOx9bgq
JGpybS5qvwWix66Lx+cyrDra2fEA2N9WNjA30UK65Rvihzr2s12YDMjGC1getX/NoCrWEF2GgTYd
1jwpcQXIXPxvsEWhGBtaVUspr4redHxTfOUZuKo2zilN+2foyAWHyp0q7nQgYX+tL0CpdJyzLXA4
ZvC0sg15HQLpT0DNsj10KjML8xMVAa9PQG7goYqikfSJjQkd49Ay60btCFfeTXcsSq24G1WqGdcy
dVEIoTUFKgErMbQ6Rtpqae4kn4eTQUyclybv7IjBjshy9ecb4ZsxPe86wc3SptNg9UwVPOqR/9cZ
0XGnyTFWlFc4uiHiwHo+Eryl/ejamhjbzjsA9a2o1cBDbtZFx1tXYksZwHK9Z4yJ1IpBVckabLfq
jCokf1/D4NcfeYmx6DgVcPhmkPK7+fAtiAgmtbduNq0xy5TCIdlB6VniQispCRIUOTvfRw4Ut+B0
MgMd8G1Y1VQEoJIc/9Sgx2hd4cDSUW3mva4i3kVwR/YYMnErhixfL0eRTdXlwQ4bRrVZajcYjFu0
Opg7H6NZnD06SjqTx2eBO/zwauFjnTrEMjkl8RV30beKggOIAxnz1Gt5rjK5lPUvX6Idm3yFP++/
sFjhd9E1KeYIYjwTEbyrxv7vlb0QKTDijMkCKWfKEgy7N8mCAGBNX7QA8k7imhf2S30a26CeB8cb
Jl6panNGdTdjbEcx1VhKC0uxn6ZQf3jXH9YmKDOYHp5HdVeIS6lei4KCeLxSjffXp/9WA7n9gJ5q
MS4ezkOFVD+3aNjKMGvT0I/wOXcbCSf+VApUKNrqQOkoT14ZXdflgY+VUJWEnQEG2m+XoBlZeP/x
r4o2P4mRhBcvkDw8qcz7PmjrZtQPw3MPMvvrmKrFlx/7Ra5RKuxGij9sGQNy/RzkfpopYT/mMoDr
R3OuJGN9bBT2+LRpOaX0Iy43W0WbIfGUsdFrIgIkfW05nakFSCqcHWMYYZNCeBbN5y0+HkH3p7uf
SkOVqlcJwWC+/Anhy56HpPHsi8u/YACcEQeq2eZduxoMsEa02QCvB3wIpcA78vHS+78TmalHcVA9
onCoD5wydTkgBHnX07FPENrl+VU+qSknrzNSERvqBH1x6OdfBjI4EA3bxXzAYv0E1F52CbEK1MNe
N9Ehb7pU
`protect end_protected
