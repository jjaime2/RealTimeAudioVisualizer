��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊�l*��K����C.J�_/w�SE���#V�����0�$��_J_2V�4R5��7��������T��ʵ�!��1��cx��UQ���j��*ω\s7�'��5-�@&�:8�k��̑���,����%���C��X(8tU�p}SJ�M�	n�7"$��fH��T��@�,�J���#-I)�)B�REa�O��p�4�5y������Par��N� �|�A��c�F����\�k�>���w9&�`�B-%��B���ƫj�N�
�IS7��%�sB�S$Kl��3P��D:u�����}�[�=��D#����ۯt��-M���3���X1�	��A
�6���5�?�|����t�&g!�Oƹ��¢�K��a�a�<�&��g��R�ƽ�(��4r�>tB�nu���0+#%��G{�!E�`ؔ�ۤxl�~������!"��K�|zȬ��3E#���@�R6�aW��>Z��GN����+#��k��Ky�}�x�-�;I�h[�E�	4C(�e��`U��)�߼Z�n`�c��R8��� �X�)}��x��(�kǻ 9�uت�������WƄ��iZ����4G�����t�&��3��Z�{tl߽\F�B&�%'t)z��V�U�Dx�6=�w���Binaa D�v���g�5��K������d=�Je�2"�8�a�K��]1��UE�o�c9�Ýeu��'|��j�:��R�~"�_����U/ٛ�Ĭ�6�E���i� ��]2.t�↪W��<w$�2i�?��Զ9�9 ����ay��@��y���6����}�<��{�=����H[��E��0e�j� I_I�������y�B��H�ٺ����ֺ��Me��u�;�j���ڑu��>��ђˏP(t#a��`t���>�7�eSńO�W���.���N+ j����A$�QK0R3F�G[Xr2��4��E�u����Qa�v�lJ�3�Q�G�x�P���t�m'3$ͻ� ���q��s�D��"��]���{�"��%h0ޙ���6pV�:�y ��5�ͤ���&_�>z a
��0�r�>3�V׏P�E���7�|�)�$�Bp�m)�����R닸�`�\;�DwG)����ː���2����ve�X��y]%�fl5N?�Ԋ������T���M��J�7@q]u�~X�1G�����:�ɧ,�9g�SDr�&�~�Ɖ~����1��s�K�xͦ�@�4r�H�'�+1��#�X)�d��_��Z��Y(��u�y9v�>O����w�r����F3�Gq K ���.�4 d�p(�.Q�O=��3E�vl�q�*�v�r�J	�B׌Rg�`�q�q�	֓Rf�^�VΤ�^z�����������5�?��� �1���*9=�4~��
sk�f�u�rb�=�`y]��ۘ�ۼ �Ǉ�K��g�z�"Q3䯟`j?�u��?�&�)#ąt)�6D�0m�v�aD��f��X?_}��T����\���BJ��H�,%��wx�[��E�H��L�1�^	)�$lS���O��e£�`
�����Us�[��l!)X	�-뿃jE?j�/}%����=e�#Pi��$K'jaꉕ�%Km��/���q��v,s�x�tyB-"Q,*��,%bF�k󣽅.Gζ��<G� G�X��e����,_���P|-nr�p�	nq��_�q7��&v�X�FZ9�=Z�uMX�-q�lo�0�\��̠�Wf$8,-�6�����$�Q��%Z��4ùa�$�S\��!�13� ��h���_b���b>G�aP��G�3F���紌E�^RW�H鷾D�P- �^?Y
����>���o��"�����Ik}p�'���*���u�E^_d�����:y��e��K�����N�'�A�	9'�c��C�Ɵ��u,��H(.W-��	���%��n�͗����09� �	�4��)��F ��,\D^�`�l3����unR�/��-�	<P����B	"��/n�����(�2��)�'�u���_����P%/���(v�P3J�0ѿ�?P�`Jo����*r�5�[,X�V�.ޯ\U~XS����'f��>�n�rJÃjk��w��X �a��;�/P��#e2;��U��.�\5u��a֑8�~-$�q䷖�$1�#�N%B�:�@G���;���LVaF��6���&*\�j�⭊ĕҒgN�UdfJ1&��{��!v���[�|;#�;�Ac�vP�Q'�N;��8uEE�ʭȫ��#^s.�_0����xK��n])8nGq��zM=�.A^B��9��ꃚ�����:�l�q���m��4��<f�Nj7; ��CM^W+l�R�d���r������>+ggW̥����r
-� �휵�*i}����~f���D!����Sщ��i�z��6�&,��ؼl)r��~�f��5���l(B� ����:�3��=F�$9��d�(Ǣ˔�^҂t	.�Mr^Ozw<w9ԏ]O�<-˖��<�d�@M���d���d=d�%�.fq_S]�n^u�������a;�!xג�nTR^9 ud]�U�W*�T'�`,���P� ����Რ0����(�Tߋ���qyb��d%�JG�����wV�~`%�&���9H��6E)���:ۮ5��p	v��QCb���+�'��i�����x�����]�c��ݲx�P��P�K��q���ϐ�%S� YL�_c^��0 �����p`�Т���/E;2�%�3�I������X�@�uObg�e�0�������6�^V,V���Z� b�E[�n�8�K�C��Q$��O0҉�bF�P�#����������N0&	��{9j%{o�2�%��}�[��ЩTm���w#XM�eu������ 	���".�� H�i��>e��<mjD?���"a���6 ��tƎ�
�bCf�nFX;L�*�C�rr�b��шH�s����X�iV�<D�K	g<�z�}I�� ��K����oZr��4���;�B��jw�EU��aS����Lî$c^C��?�h8���k�\�Fj]Lq����4�|�QP�K,��mb�9ƪ�������<9�[)�=��3��c���:�3rjõ��@�O�S7)��k|O�g�f�����43$St�8��J,� ���2��N��2��a�aJ�FA�����������E�:�腑E���|��c�!�N?K��ʫ�uL.�'��*{h�� 3אK�b�޴j�(��YK�Knϔ��F}G�ɀ+�R���eԼu�u�"�Zb��3���Dϲ�1���Y�ĚE�,(Xd)�U0�DN+q�Z �h�W��J���UOZ������dw��őh�J��H�'�!��$��8-.�8�Ӂ~�?D�2���A�9"�\Eql�OS��	3�����/��x*�C�5nIm�ܔ� ��x��(��|u�)(�=��>�4���#�@x��f6J뇐��\&�K��eQ�bW���H�r�n�`@At��휞��KR�`��F�.��4�ҏ�oǕQ���X���C��j4����+� �����QSMl�Π�b��ׂ�zy�aX�=�]�� ���!J�����8<wFV����b�8�S���D���z8�C���'b:|5����I"jy<+JRn���y�~@�ю^�4Ø�ҤK<?��m��^�'T|ܹ�G�
�pUE&J����+A&�]בF�q�}5�]ǭ�`t�z<���M�GT=@�kS�"!j�Q��
)>GL]�"D����m!]��72*�>�ViTnyԺڅ���V��1F�W��)2��W�ݢ�-��a�
D.�m�S�
�c����׆������_N��
+�K� �- ��=G��N�U�ϥ�wg�h�v4fK]��pd�i?�C�5���l�q:P� ��"���@ېG���*)ѡJ� �	���5�&�v7K?�Ɵ�L�������x�w��=r�
�p�<�/���$�K��
�im�-���8T-8�q�����ٷ3-+@��1i�^ؽ�a���k�Y��U|ܙ sX��0U���W�Z��d�)(��~$����������[�6�=&�D&�����TrM�<yw��%����t�J���F��]����(�
b�]A���e�s�bf��H�/$��� �7(u�S�'	�u*i��&�^5P�rn���s���4���*Z�zJ�����YѣG [..�e¯G�C��t�_��)��N�wwK��|#D������/1�*}.'/p�v���'3���hw�x�q�n1wl��aG3v]�D/>���l]Y>3�I܉"�}�z�l2���m���+�}c-�ҳD�3Y�!���sV9�xM�ٿ��������:n߯J������O���H�j�����a0�q_A�]�NV6Fm�!/+3���,��*�Y]��0���_=��	MZ{ �g&"����aFs�C�f�k?b� pZNW�m��A�c�{,����9�׎#�`��~�U�o�>�3���tv>T�(m���J
�>���ht�0=�]�'��T��
i�]#*׽������E����4���e�~��o��i���H٥�
a��YOeK̈́|����`��,���u3:�#"W&��Y��-���M#�pR��-D�Ψ��՗�T�7��-F F��[2|��o"�ѣ	�}����2��>wbq��K��9ɜK{G�b9��Z�3%3�m���]a�N �3����=��s�w�x�4��1Bϑ���Uox�a$"ki+p��j��T��;��}��I�7koB)^|���lL�h>EVS�`v۟�G��p�4�G[�����A��>>SRtt�Įҭ�<]�����L���8��p!3|�u
el�����!"��V\"�}ԚQ�y�:�*�nޞ�H���>�v
�y
���L�}w/��o�@j�=־��pPZ{+s_л<�k�C
�'��Y��Jw�с�Y�7cM����(߆��0֬"d`��$�c�]O�����������P��(_���&iq|�6$��c7k�@���h3��^�3����9&�b朠�gӧ�ޯ#mķ�D��Wk���6
�!�/4k�Y�8]B0+��h������s˸�kE4ɉ��՛hs[Q]=ڥ^��>�k�̥ՙD9~��/�ٖ���i$�����Ħ,`����w{�TkB��8�ș`"p����m�4�an�$��ا�0˳����1����8�>!���ܓ7���p�c,�ų�����L��c���hm[�'|(9;ii�QW�Ɓ~����������Z�Sfu=���A�`C�d����?�`��-�V�߀���ŏ�4VZEe�B�\��!oe����r���[�X:�q�L��W�A�3�v/D��u�W��C�8$�ʵ���'wdt�q.�O@�2����Y�ŝ�����"a3���ˌ���p���J�w4!0��=w�>���mc*�O��R�4bQ�_�}%�ƛ��Ջ�\��b�N�jt����M�\6*{�ۖ./�k�o�`w�i�A.o ��i�@�_��0w��`Ǘ�4�ޖ9�����dWcOL%خL�6Ym��ux���N;C!UĴ�l������{WE�fhB�|�@���[Mp1!��������a���~41H�<��0��� ��J�.
!Il���TP(>��MP�Z��ظ��
�p�*�W���G��=��w�T]�žS'�6���,UrX�|�k�}�z-],����t�����6W�	�`�u��C����1�,��wϺ�+�����ص�1
>��( ˥��dQU��u��܏.�{y��d��m�D�G���Whb�Z	{��nVo�>"���]�w��	��(����<eYM�퉩R��>d�Q���< ~�׵ &�m%��<�Y!�l0��Tw68.��hI�,]WE��νi���ј����ؼ�.�������t7Mػ�c��T�4i:+�5Z��lo�\9Z�d��۱_T�3�������{������ȋ�:��$T^�d�-P��\�\���o��*>Л< oh�9���;Bg3����F6a��G�o!y0w������άth��y����?^�˕�}I����	�s�D0%��-�n1�S���l����1�az�g�U�ǒP9l��12���qU7�����ix���Nt��g}��+���[<p��U���j������.pJ��cDkY�C��y՚�e;�(�h5���Q$�����j�Z0m(�~�O���f���l!����cH����y�*@��O���<��yt0]�����-.QWs���G1s�f�C�H��2&B����R����A�s�cd_u^�[�G59
4+��/�#�D�a#�FK�:3L�f�I����:�It���;H�����`E�	�	�*�vs������YO�� ��s����a|����nٛP~Ǫ��F�s���uy�
��4p�TtJ�aWLg�%�̇�(`� �� Q�$d� BA�e�ben�hv�ai[�\D+]|��W�҃k�I/�0~�?�������� ��x�IV�u�ֱ�؇�24�ҥ�'��,)��\*��J�S��#�x��[�
��K����ԁX�����N���Z6�[�9�T��1A!�/���E.d�@\�O�[B#��2	��_i9w�ϥ4�b��1v,�O�ej|{��U��?�_K���#mUO��2�ݟ3�ed��oMX��!�Pt(e-�J4�\J��� "~�;��uf�}M�,o�,o<
�~�������KF�D<�s:����Oݺ_E*�tL��v����ʶ
w�,# ޱ�@�#0��Dyw����r�ۍ۴�q鼺��Hzt��9���W��e_��Rl�n�\�p��Ğ�H��i��L@���T�!� +�NԷ�1��׎��H�$��ũ�@��o��Nm�i!�r[ r_�X$r���A;�aV�����2��������[�"<���aO��P�	�-/�瀿��Q �ɮ,���(n��*��W��D�U�<��G)ƀPϿ�-�#��U������*u�x<cG���S�/��6&i���<���Z ������s)Ҫ�K���s6 �4�D���T�_�����|�P�S�>��4��A��������kM{�%۷��E����Z����}a�Ȟl���!����5�]P4y�i����H71�E����ۅ �M�A@�[%T:�D������n T��pr�F��>�k�p���q��ұiP�E�~��9�f9�lq �$e��4�|H<�b�Q�6�����_�7"l�"`�p�c�kЬ�%͆\5���B�#Y�#gX�y�*~����"Q�>��l��*�~��  �-�Fc�b�̡c`�����u�xc>G�r���J��[�Av�r��Jb�����ʂ57�'fڃ�3r��̲�����t�Nf]�,>ฒ@�������sG=��>$�i�5�^s�4��m-����Q��!�&@���(9w�%6w|��g\���# �9�X�,Q."��3�gy>ǐ戇�41��b2i��,��<� l*t���鐋 ��A��U b�yEp�����W̮QI����������?>D�[��%٤��T �g�cNe�})�Hq8|RI$}]+��~���;l�ɲ�HH(�t�N�()�ȧ�I���%�Z5V� vb�g��BI5,���>:��ƠS( �n��_��v�$������BB��	��~��L���t�0I�R��;�N���E��۹�`�`8��*%�,���Ѫ:~礿G�ؠ��?g�K��'�uȸi6������(�.fK�:�hMi�߮�����*��}���հ�{E�����0xH�^L�0wPZ@�S�w��dn=��=���5��G� 滦�E�s�2�h�T�$���'��8�5VX��)o0q��y�S�?��0����Ko�a��@�ڏkΨ��>Ož��s�H�Wx�F<�.)�޲e�G�Ew��	�[t��b'�9#mC�_���8�z���L�uഏ�P1�*kƸq~���YZ��_�R�sxX�KĮ�a��_��7��144>D��b�6��S���#e]���r��89Xk�}�-�P�>CW`��3$DT�e���ۋ��S�.H�L�� �K4J�s1?ņF�,Er�SI(e�&���?�L	~2�Y���$��5�79�}�b؀�����Χ0���\ղqП��fC�(��
6l�.֪*���G��D�(�j��#3B<��8B�+��s()������&�5Z(��������1p�0B��8٬�p��B	�Hګ��J�}���"^W��?ns���=�����K��ޞJ�/ �l\�����<��Q4X��
j�P*5���N�M��Iy���Mg+��qyȢw��dN�R���!/�h�ͺXU(}���ʢ��.�E;��8Bem��ZL�j)�%y���/�_Y�b��3���Y�SR��)}�anP�>����u�y��"���5���'��bG�P�j;���Zq�*�E��W�D�'�����d!e�(Q�G֭f��&!W�Z�葔O,���@����(}�vck�M��\�"�'7l� Gw�n����!�hy[�1��!�r��`����8ߤYH��d��gv����t?v\�����]�F+
<W������Xx�b�PiJIm�_m3��Ї�6��x�[��}�+���b���r���O6��K5x��\���٬eTJI�Lʩq��E�jo�-��~���d2%s��O�N;%���f+�o6�l��}u��^5�����Ի�E��o	��\ŉڑ^-0����6j	��Z5y��g�	���g+����ž(����ѐ�:Xr~9>�D!O,3��6�)m?y�����Ǽ�p��l��K}�.��RIe�Lr/�?�J�%FHAFXº��ͭ��o\/�e�j|���笍v��z_⤬Pr$}क���)��`|��P䫺�������{ ����Q�EJ��`�Śi��l#���YDFu#F��B���G��λ��#��be��Ȟ<�[;2���G�#/�ה}���1�
����5� 	�#�X�����?Lި�P��k���+察��	ҿf$aO� |$ݩ���HH��ƚjar��7��
u�]	��U.E�l������E�o��)��0!�Dgv���0f$���lɶ��$�@3��\w���$��~�Y~e��VQ��GS��@2���k,~f�Zg�ਭ�|���{�72��5Ed�Z��[�;M�{x�;�6Ӱ��e9�i�J�n��2D��ˉ;��3���������O�Xf
jSKL�� ��x���	FɊ;y�+�E�2�T���L%Y����Od�<��Q��J+A*��D�ЛHJ�s!���:�^6���<�����N��y���$�i�k�.��gpI�3��o���X.�����C����U"?F\[~�p�8�dqɃ�./�RG������\�(�He�
4�Z�������>I�I\�A�$"c�q���Z�U��h^� )�CN����U�6�*��2!ԭ����Cf�l;@�����LF�V���_t�X�5�tZh�2�Z��B\C�1k��W��?�[i�Y	�'	&X6kv��2�;��z�m=2X��	S"�ʦ���H����R�AOk��qڸO���ᫎ���T�II�!�4���xJ@Hf�8\����3�Km�L#�Yi�� �Q��U��d�Ў�jy��F��~,6&\���W������l��}���"��7t�*zj�ٽ�|{�j6��d�u`N{���y�L���7'贡g�����ȣ_�~�Հ�EQ���~���qJ�SU�T(�ݖ��\_���t[��JD�pϫ%ђ2�j��A&�j��u�C�B� �`F�I*^���׻|��b��T��$�? ta}�d���K��p��p��4��r��.8��6���\i{�g�o��&�`hW�q���������-�
8�������Et5���I����n	Ιt~k�Dcֱw�.ˎ������&�.��䨹9�̅�ì3���W�3c*��
fu�C9L�}��q+?�}9�:�i�r�"i�t��EBR$Y�6j��/��%�$����j�Q�d�^��𽅞�>��_�κ��� ,�\g@|��d&h�xm�tVP�h�Ҏ�yD!�����GY����n�:������0���~H!���z��My?�]��"^J��	���v	f�f�F �$���e��j��u�l���m���Z�� ��w��ir>Q����;�^$�78W@��>䫏N�����ỲBNJ�i���`��O,�=Wy��rfBiz3uڷo��[��_�_��3\�*J�B"P��V!��ja����*`�3$�4~C�Nc8�(GUn'�������|�bN���3�[p���3Eu-�5�X&�L�q7�������,Yml53ʚ{��OE����� \��tDB�w��NQ_#�Y��H�oW���I3��gU	��Қ|ʭ I�[�L�xF�������3�tg��=�gK~ĳ {c>���4�C�q���-n���C�(/MKԣ�U���,��
�]E�lb�o	�(X���nW�kb�A���,�١h7�t3��_Z��j6�r��+���/좑��|�A�� ���|f�$�Q��-�Wh���g�v���n�M�k��7y1����	A�ޫ�c0�ᒯ�|���m�}����ȡmS�;�|�v#�^g�G9�I�S��P�5��ԭn}��`6�-/����gӂx���}=I4��6{>`��'I�4� ~���=ױ ?�nec����A��LH�_��_�^68����d�v��1;&w_���֭�ƾ-e�$ ��%״fz�枆��l�A�x���o���W���Ǩry�vM�$���ѣ?���F��l����(}>�"sM	;���z�Z:���ud��XM�q�����|1�cުo�Iz���3l�\ؑZ\�p�U����?)�ẹP��m��+�\u*�%�G�b6�"�X9���Z���e�oD�}]����@�^	��$�D.�EU�>Y�}����_��&�F��CjV�>}��i��fE����Ю߈�F3�����BE�U��5L��˝	�Ôu��%�_�Mx2,g'���k��{�h�lJ��詁T9��2<����`��=��<��rJm������D������$}U�M	�4L�)V&j0
=��T��$��
�H���=Xg���<���G��T�R2������M0UD�����$�4��>�*R�	v���~�Y�^Ҥ�b�"@��&�t��D�]��R��d\��扤Ŭ������2Ȏ�,����B����kų��8��:�i�o�u6�f#�g}�4'�Z|G{��P�ƙB+�V ���Za� ��T+��G��^x�,�_˾ʾ��_� �W�a�ޅ�\�1�XY�4<�ir�j�F@�jt>-m�vP�}��G�0���&�|�q��%ح�tG�����]l�9:xT�W�3��4L6�q��F�]u"����~dw4���rV�T�Gf��G:�ٜeZ���e��բG(�`R!V@��3z觯@��7��q����� tيX���י����IX����i��S��IQ���T���G#��ƍZn�c�݌Anצ����R[�9� ���ĺ�e��l�~�T����ă��csE�NA�"R�7��7=a|�B$Po{!�V���K	��Ǚ�3�尻X1P�*�v�4+�(vZ���1��c���1@���$��2��GH B�z-�I�O �q��@:x�I9t@��c_}b�fL|m
��\��
mP��;����%es/�9%��	Nf��O�������X��� `TNl��~w�0�w3��Ka���LG꘧aS.qmF��:E.�b��a/^�DZk��o��ȴEC�}H�E��T�8�lbK�Z��u�
'�@���z"��\dE.�}@ʜ�	��ݖ�yȢ4�	Mkm�b4�5B]M���ثz�5.�5�=X����aZ�����q&����C��GL$��@�h�bY~'|�W�u�Z�]�i�'���$[#���$��CM��x�A��l����QA����d���⑟Z�q,�D8ͅ�8'�0�g�:�ڍر7z^m�M��� �h.�������)=Ѳn�˽�8�g�1�%����a�0K;���w~���Mό93�}��O��uVb���Bw�ԅ(��jP���_g��Y��U�*�r�-JMro޻*u����kl��[�	.���h�.�1bX'T�����{F�!HI4���&�a�#�$��i|CY�FF��_�V@��^��P�.=Ӌ�D鿩�J������]��J���i;����耂�<�I�_鿮ٸ=@7��T@�i�Nb���sά����]��>�Jb��S���*�5����b,R(�J��j�����jW�ar�\vU�斔��>�B�{@,?pW&|F��d m�����_0I����\������/��,�E��`�oln���V�D;-����웅�l�������k=���}aˤ	G��!�$�۝T<h�k�y8�� 0�6�^�ul��a���H2~�v����#0В��t	}�W���.����}��Z�$��9*�4�|kPoZ���l�^����hm�1�LL��w����q�pU'W�׬�T�ėu���1V��/	��;���s3����u�x�mj�K��y|�����{�c�a?;'���o�J���
���|.����9����(���n�%�N�Pv�U��wl��q�F�^Xd���\��b�W�Y��U2��u	������`�������M/�I��3����v��"�M1m�u�"v�Yf1X�hJ�ɹ�*�۞�uX�����M-1�6��� �����?�,���d���)*������d�[U�������j�i�`zu��1f)�䋜���XO��Y�(�j)6�F�Mh@�7fðk,�����8���r�T\v��<�*p����/�����`��ϋ�.:��_!{������w�4{M�I��\��Ll�F�2�m�t9T����\BJL�k��JM�f���4|��׋~��r�=6��jY׻y�G�P�M���˱��
�&K���b��Ѻ���� �B�^��ʨ��k38R�ͥs~��2vKܦ�\�=���x����Mk��<�
'�鴃-'E��j$�����mU#'�0{�s�VG���.k���y�.3�@)�<,��'�o��V�ʪ��0T8�����ޱEi��t����i������Ь?h�g ������b?9w�FW�Od�F����R%���ܮ
e+�.է#p�ۀ҂�z��r������(���\����Z� �z����I�y�!p���������#���O�ZUu�}Qs�E����<��XZ尀���:�0>�i):����zu�BL.���;�]OI�P�m���i�O����]�'�=v�9o� �E%���--N�q�<�<��j<�RV.U�i�u�>����M��Ō�s���Z�����1F��onC�pO��#@�F�d$� R��2.��Z���
�N͙sd�f(B�*�?����-鄖���pB�H1p��b��7�R��;�������vK�~��X+y�����<;ot���eK��J>'����޺L�΂oP��^�X(O�h ��	���]t�+���B
��K���i�q�᯾��l m2�":ޞ{�m�ٴp��&oO��.G�l7ە�8��Qcz��q��8�����jb�w��X��<[��1����eH]�M!�M���
v+(\y�Uѹ��b�`�v��X�>��|ԃ�b�� (JH�q��G������nfd�N섉���q dщKh>�����8��4�uA�h���Ō�W�Pd�M��`dl(L��dU���� GjM�"�&���]��=�k[_.y��@��	��WN�������'l4��6��a���V�~҉�E����i��b�ϛ���S��1��^Q혋��+�:J	/��)�J��0�bSb1)�RD�5�o��aܬ3]Z9�=�q��:��;={���˻+u�ɼ���55��ۦ��d`=O�6�H��{���h�K���y�m��@���h�/�����~8#�UZ��B����S�u����$_��!Z�=�)�������`� [��J-��&�_2��c/b2KKVO!�a�`�$V������E�8��iO� i�����,�D���&t�p!h�$���g��jmPr"����]����>D�Xk׵�
�O�5�I���}���?H^�ľߋb ����^�W?�h���jU��hzM9���I�Q�����W)g�Y�B���0����&�vy\R����=v��w���8ҊjE"��g���~�\���H��j�POL���Z��{����B����ԣp�j�O�VB?���2��%t�-�r(R�~������ �_��@	&����!�d�`��';� h�ıT��amP��K�i�#Hc[�*��w(&�H�D�S�XD���Z�_�LƏ���|���;L�I�u0�{Gfo�pR1"&�f��9��J�c�P+ix�p���>���oy�z�\ ��J�W���q����ѹm����F�^˓�F���a�k*�8$Q\QX�$�/d�?�1�������Dr�&A1SRz��N�eB�^�5���,q3N��`�)� �}���TЍ���RoY�/�,��f�v'��ih��F*�h���a��nr5y�fO �$�h��EF9��Zb������m�V*�J�k�|��.('�"g;0���cd�yc��B��B�rk&`�wn�������	6��Ό~�Y��6�Z ��W�>UUX�	�SYc,o�u�nU���&�Z'�Ae���FȖ�0=��+�ؽA�:?�[����f-�3:5���j𺷕t,vc�o�C��u=�_i[I���=����]�.�i5(k���V�Jgg�� �N~�7;��BW}�t�T�	�g�Ō� �0�C�k��&.e_��T��B�̎�&G{�Lg��\���M�(��}������,G�m�}T`��]%6x���?�A,s���Ui�/y��!5��C�a�����m��0�>���G�qe��<��LV;�¹��s�!�f�|,�@�a��,]5u>K.Zp�z4E��!pN)�v~]��=�@G��϶�fZ�k�4,m�Ȭq`8�31b�O�ő 
5�t�0A�91��^��y�k���G{�V(Q_XHC����7+
���;�]�o��������˟��1n$̐��� ��I��WGe[�����e2τ煜�4vW҄ 1�!�+�g��@����������9]�f݄6�j��-n��
�[��0�"�l����ycQOK���J���*m��~y=��?�V�1�T)?��9�[K�,�w>z��B��{��Y���ʱ1��<X`!0���zt�	��̈́��m*�. �ݕba�5:�?%dR�������G��d�<��nfE�"�L4M ^�ld�dG3��0@���1�������3���[YFY\X|���i����ZcŇ�U�w�ٍ�%Ya��S��&[�|�Y=!J� �X*L0g](�ѱ3�ʾ���/��{�X�g�AQ�{X�:\D���T��3t�3�����%�TC���]GJb%:��)!����a@	|�D@'lF��,��GM�4ڎHd/I��?Z�ib��6a��H�GA����{��N:]�n���n�q�&_ ��`��tu E�B@;�5��нJ��ˀ���c�@S�N���0��86����rΫm��*jͥK�G�U*�u�b����?��"n�`����@��e!x�-~�/���tWy�(ddB]I.dz�(����h��sr���p�ύ��9˩�f�k;��#F�f��p8Q��'\�~1���-���ɟ��t�f��1k�ќ"zs�S�>�lC�0K?��&��7�̓�4o_�bv�4�k��x� ��jq����@M`�0s(�	q��Gߜ��i�)��8p<4�y��¥:4�);c�#9�ų;M\+�<9�
��-�pz��V���%^Y����r�����x� 
i����UЖ����n*�m榜�:�Pǳ�O9�̼��3���*�j�9	DV��01:ۯ<�6���z' �4X��x���1@1}�C��mu-æ��ՙɪ@MP?O�N��5��u�X�Wm�~J��w=��V*��ހF�֗P��G-GL3*�q9=��<�(�d�'��h�{9{�~�}��E�.Ȯ�fg�����.QN�D��i�KԬ�(��#)��3|��z�֜+9S�5��]*֊Ǆ����z�Ϯ_d>��&����:�w?.@d��x!tw�v�Г阛{5e���� S�*�&�6�lYA`>�5� .�RyKKH�%'��O��:�ڗ^��)EMY�s��G�UK�2����79��%R*V�z�Z�x��T��̠d���`Ψ�cQ/���k�O�~���U5��C.)��`1�y&z΋`��wV��M�߇�����s�)���{R���[s��Z�/8���n�?�r!�W�.;��Ct�Cށ�� Q͑��S�`w��t�@	����8@!�1-�R���ԧ���I�L#�
�mZ�,��<[^Y%l����l��!0���Nצ0�l�� !���0���F�;���,�t�H�{nP�j��X��'(l��gԇ��Y�.�J��bK������qK�(�5KG$
u��;��z�H���'�X���q6�h��=�÷�3iY��]���],�%�U�S`J3B���'M��){@����klr'��{��mm�Ա����8DǠ�Q*+�_��7��(W���,��׹��P[�0�">�Q�$�u��3���ɤk��X����y��4��U��o|Ą�|�:��n��,&�Ɉ�뤟X|,����?����s�Q���>��������S{k=v�r�e߇�[J�mM�h�<�OŮ���2Fr/����� �K�'�h��UJ�^��*m�Z���%Z8�̉�q<���f�̔��gG��|Ol�{x5�)�4��}�ɻX���iQ��x_����7���Z���4w
��ބm��=5�`2xG]?o�d��GE��*��-;�&�d|X�'���*i��Ȓd��aycQln��׃Ӏ�s�����̴6�xyɛ��Bi�Sp,�rܲ .*h��(y��k�
Oϕ�+" ��@��g��T�^���6-�Wr��&�
��ओZ��媬I�@R�����Y�Z��#d����Ȉx>}��3(�0���4�H�3L�1�����:��W�|�e��R=���.ʇ.~X�os.�������h�iI���^eF-������ce��+gu�'�kP�X��.v���"����1��}*oBcs�ۊ���@�??�\4�{��� ci��h�ka�T�_O���-��]�n�*/�E*�A�Z<����	5�I[p�K�x|�d�4��:��/H�(��g�qj':Y11��Eՠ,����xu�a��,�dKv}|t�����ơ
s�w�ϋhs�Ua���D<�t�,��Z���ppa�'��f�p��;�(]�Q��Ƙ�h{�ߞU��G�6����bh�'5�{E��?k�9�-\��詝}�s��P��l�]�A�٧�ۑ){��e8R���tݩG���^�&f� ��Tȟ�5�0׾�p�*:�!�/(��O��y��a�G������v
L��S����.�J�Ĳ�eU���s��G��%������H��h��4�Т��LF�v�h��`@XO�N�"� e�0�-�?j]f(L;�*'�y%tv'c�c��?�HF(��^�����ߥͦ(b�[�[�j�dl����} " 벜=�{B��ȴ�r��O�͍�>�j�y8���v��V�H���k)YuL	_釒���h'��(}=/|̇��J�kb���M֒�����6J�y�gN,xAf�z�$@?=����w������ø�\Hl7����0<ǐ�E���6#���X�2o\�w��UBT��61ޏ���(��!�lU���qCI���dE*x��M[�"�
��2?D�qZ1��ϳŁ8@͢�_t�ć� ���o��_ݫ��e0�)���� wR�A��?4� �q�A�mf�Nd3!��1������%�ݷ|9uc�>o:�W&l�E��C��K�;*�;���H�˗+�l�������n!u�p�s�6w���y�4C��HewC=O��Pyr��?�L����& W~}	uDح����6~[�@S���*�n�n�Z�4������XZ���=5��fS�����_�R��CX *|��}�?��/�s�Lw��+8��C��C���C�kUP~�E�����%�x{��^����,D���2�ɐ������w�����t)Ⱦ���R?�W2}���LД\�6����4Ggީ�^(�_�W��[C4B]��_�[�&����D%`&�o�����4�6�駡{�kAG�.
�)p��RŇ�z=�;ɣ}:G��0�wX��<Q�� /Y��ZZZ��W�Y�CY:��A�̗��j�O^��6<�c���(�`W�w�)��+.n:2?4WH��x�
��U�t�6��N�m�UB�')�r�h�*���DL[]��Hs#�gd����gg�^���R+��⫎�96>��	������i�|5y:E�\�;�YP�P� $���O(�p���ڏ=H����/b�QRC�)	�$�˟��R	���;���G�I����p¯�/�(���0*��q&���/�	��|el�L<�ųб��G	��(&4���u�@�jȫ���`v��m���_�f�n��Q�o�fwl[u��!c[�@�kҡ���#]��5q9���:��f)�)�Bǒ��@bǒ�M��ԡp���ʴ<@)��]��d��ܕ��p�[����
�b./F�xw6�T��u��X�G8}D$+Ed/�H>���]�����2��0�w�/��0�i��qj���wC�:=_�D�r��<~n�0�pi��z}R�=L���Y������Y�!v��a�hP�~��֡X�����u�{�*
�a�I�.��l�K�	�Q�<��ǢR�c�cvgL&ף0��� �E[��� 8�
}��KW1H�u�:-w���Nd��p�ĺ�0GG�E�oiӓ�#�y�n`�ulgU@�k�jR��,�<`1��#�oۄ�yaC�;�RR��&��⦎q�(��0�"�vZs^m�Sx�����Y���Mn�$��C�4i#|5�h�
y��}[��\a ���C��D�.p�mv�๝ʂ0k���J�� �([��8�p
�9�(��m��ؒ�������RU\i�5���b-�/>�L!u�'HO��u���Cǖ���؇^��-�H9��#�H���f�&(�V,��Z�f�!"�w���VO���S���M�J6̙4��,�E3�u$�ˏ�9��PD4��V�.�E�O���z�=$?Η̞Q�eJ��0��`�M��RڴI����S���ؒDk���`�|ǭ�l��j�-	�\X��J�\����U�bFwT9lB	�)������"�(2&k��Z���&mrM��Y�5*?=Yl8�i�
��c�F�Cd"��3�����x���f��V��>���f :�X��'�?�u���,w��+`�m0�aA�v�%?�0��Į��0$��$c��_�z��I{t��Ed~�1�i����OҔ/�&��_�
�i��	S_�xL�Z�,�&0�4����=�hTC׺�byo��n��s!rT�|zޝ�؏!n{US�~t@�qgU�lڕ� ��µ9{��J���:z�*�1Z����v9�XB`Ć�_�߯o��5�����n�K᷃����L���v�/adAh��EZ0~|n�Ⱦ`c�磃�<��tXw�2n��p�,��K	ʑD�pB��ֽ�b������Ȩgv���a���:(�<L�X���]e���NH�Y�� C)�) ց�w<Y%m,|�,�Cg	CN!���ĕUr0��)7F�#fK$��E���rm���4�Q~�ɳ�v^�9��Ȟ~���2�:	�����	�((w�XwIk��{�'}�W�LE�nHp�PĴAk<uv2�az)֝���QkA�X%
��:�}����B'�X;xF�8@�Ov�>T�<U�ʁ���k���U��si����?Љ�Z�&[����T����T�@�h	>߁c@?=OŖv8�zn4�����c)�c7"��l�k�A]	Ȫa(��P�̗�3-3/�H�A||C��&p��
{ =*�`4�j�,��R�2Z�{����~H������ςW�E���46xH�5�޵��K�4�\�Me�AP��+�/�0� ��^��#�Ege�<^[�"SF<��py�2����أT���Ɩ��!r�P�X2~~����.y��>�l��k�q|�Ls:�3��|�R��w}��F�����4�� *�0�uj����#��p/i��҈U�H�^�x�r֖ ��qL�`�[*'`������ �d�������vy��@LU�������<c�d�b��}/)p�$�'	��4�$��4f�eڷNlÆ��It.�B��G46�w|����B���z��C?�{�x:!e�-c�(ea�U�����W��ib<����@e�6�e��H.!<P!v���].95<�NS'��y�o��o�pm��r�1���%'E_Y$ٲ\j Z���sIȈ����*�k����LO�/;g��O��Plё����x(�E�;�(UEX78��^.יI�r#�����e�DG@�p�V4L�?���	�}������t	U�JR��o�,�(;���{��Ĥ/X�ǎv��&��QA�;,8���%����qԝ����6�* ��T�9X�  |qЫ���?낀f�n�Xid���56Z�@J� D^�D}�S��ybƮ,1F�W��
0��TB�;b>�ѱ��W≅/~pO�E���������m��4>��+�&��������>U�]�N��I�+�$�RM�&���am�X-u=r�kf�$�_�)7"��Hk=��ɲ;�� uEoN D�Gz������z Js#1��^��A�4�s��1���^�n�zW��f�P�r��&��O��i��O}��3�~ʐw��3.^.XX�kN�,T�q�g}�xGV�y4�͆�
�N����Ӳ�m�����ob�/�&��h+`!.�T��)Q����q&AR�tx�<Y��1e��ǲbs�E��w�q3V%l%���^�e4�2Nwx!V�k��*�E-Uq�0�61��Ǟ��q.qIˤlO�<F`=�������ۂ��)2���ұo�j�\�d^8ת�E�'�R�s&Vld�U�Đs�[M���Z�mE�=ih��N���H�7��5:w���v�*�����d��Xli�"·0)�?5g�S�GU�n�m��P	��"����.�����?�NJSd8$�����U�3��;ٶ9%o5�x�!` �F�������� X�0k��eTq��VL,XH�z&)���V	�|5����:�I:���=�����b8q�A8j�a�����͹��)�qΒ^l�4�3�R~;#L˷��,.Ԥ�0��1�_2R@��UVߠ�٪xLvod1��CV�0}w�6���pN`	�΄Z�קJ����T�U�^����y�i�|�9���fz�1�DHIg+�:�*?YZ Zq09��FP�N`!fxx�(�m�)�ͦ��4���@nO��\��g$O�ϹTI��2��V~��6%ĴT�*�C�x;4���������m�'�#�|c��b����H�M�_�
[?��K��[59е�"u���w���g��n*='	�	��+t��o}=B$v���Ns�)��z^��v�P?�ۂ��NY�h/���X��MYE�63	<�
pۣ�>��K
�d(����v� +Y��]�I#ѨX����Kd�08���==����ۉ	:��xf�ȉ���ݎ����U��\���s�C���[�OWQCa5S�*��8�K�U����:S��6D���`�d8Ku�b_��"i������ii��X�k� V�	��u�H�x��CE��	���ֺ�vm v8z50o��8eE�P/+�������ۈ�"o�4�~��v:y���D�\�	��ܡ6��e�2]899�P����@�=!?p� ��b\���3̄�K�6=�6�"�J+-'ttV1��)�<j=,�C_��$&�L�k�c�9_q�ґ���wd��e�B�P�?yx+\E6�-�!�T��A���l���y'an[Q��|��r�񞫙3f]���[1�@�n�:/bM�D��������� ��Մ��b��z��Z�տW�,7{K���(�3>��������㜞�m��;׬8*��W�*����$Z5��|��n���
%oL��~K��D8�[�y~��Ƿ���&@�"�L�_���f���K�Z�����Λ H�{�_�i �Kt�R��3A/�M�;��8�ف�-5�3���@��;�����Ԡ`�vO��O}� ;�'���L�aj�-�k��v����"��i���"'�5~a?<vm�(䀮�n�`��i��Itr�$r~[������o�o�(��-���#)��0�G|'��>g���X�v���dI����
Q,����X��z2���0@?��9����za�M4�C�VPKiȁ�@�fU_��9��w�^y`Ǆ�4~	9�4)j����
)Q��9l��kGT�CA1�@�g곌�D��)b|Ԗ
ߍ����ڸg��iwq��@�[��IO%�K>#_Lq�LW��X�7n̋����XJ�!�`�k�Z�M���\��T3��p���E$-g.�Vqz���=�x�џ��K��lJ;�����6��7��=@��u�\�b�=�珒��(��*���Y��t�$<��[�̹B��h䗗qF�q��p��~�˝�v�/1HY���e��z���+R�H����Z��#�cᘹw.a޳�NGŮu�ݔ4�0�x���Lr��2b&/�������2޴��V� ��1�$8w�5΍P��F~�ױ"��y�[�B���p��u��h��-vv�w����؎WUt������{�f��� �C�k:E%gP}���nJfS���%�q`n�ZK�I�R��M�=�%(��t��Zv���R/h!-�:R�*گ�a�k�����l�Ss�`²BW�$�<8�ѓ��F/�2��u�D�H*uHi�0��XF��k+����|��@a�l�!<U�Z�Ȗ�����g-)Ѫz��P�Rl؍�-��\�b�[}L�h�ٺ�G=W+hN��7�_�	)��Δţ#z�p?�q⭓�bkc��F��3��$�Pԟ
������9:7���)�y^��ӑ�s�!��Aɧ��8�َ�P�"����z���Ar�5�/�:&��D�m�YQR��6У����ܑ�߃l�d�~OZ=?��i��a�(�?u������앱�\�I���M��x ��7���f��Nw݄���Fh�h*k f��Pp"�Y{l�'���t<*�h�\�G|d ��ޜ	�X�/���(�'x,	¸���)+�kSO,�рe��@·��K��0�뽔?���j
槩jN{P�JW�O��|��0�&�����R��;BQ^����U���q�E]�4JL��N�a�Ӻ��0�����`��Iv.�&ؙ�1f�ŋ�;$�p�%�1�G�ض��,I᭥8��\��B\��C�%|3[q�=<���Kk-2�tn���:���	�N�xu�EE�[�o����-��9��_��y���hP,&��O��%4���Yj�'��W)dX�����*5Q7���&u#���:ae4
�������/~�+��!͂�N�Y�k��N���
T����Y�|h����&e�r<3
#��[2��1n����Ƹ�V�~��:�}Ϳñ����Q�/�ߓy��r(�K�n�4�r�dz�7%��	OT�\��ds!Amj�!�����n+p���W`I\���~������j諩��PH��8` -8�ϓ�ɼp�k�{v �f���(i7��+��S>�w���T�-���3JP���O���7�lq7:�ꃺL����w�Dݛ�6�����#*�	=�|����l:M��aai��G����i{��!����Bl@a�7�pzJ(�xN{�������p�\��Y�K~�)ז�Se8[%$F�-�*�U�͊�|��=�-�a�@�R��5o���CN�(�u��4�kL���A;����C�g�b|��}��%�.�ʑ{������Xn�yn�-W��e����%	,�`E���hX�˯o��V8b����%ȿ��.�'^��u�|1�8���E�߷\�Mc�����\��}�hk�����u������-�am�@w�p���I{������o�9�Y��E��x�oˤ�0�#���zlc�V��gC�X+P�.[�����<_�P^���by,�Nq�ťZdu���3
�<ӘW�WZ��e�Yl��������}H4����Ę>9y(��%�c7�1jud�So)c�Dp>=���G��nG��*������R��E��0j�_�'s��Է�h��L�WA��E��-W8�!��wb3w,��96��H5�[�Ɯ]h̀���h������x�J+J�z�w5����RcY,�驤��>-HmИ8 	wUB�mp�9+?:!;�������۠ʠ�+c;�C�684P�]?��;,Й�fwf���'���!�] �5�����z%E��3�V�n��p��(�Z`������.�s:D���̰��^�7ȣ��ݱ8W��5����	��d�y-+bZ=s��p�H���Ot8v�-���O	�c^���W�aW��t�F�d��d�?����	nഥ�@o>���}�bt�.�/�S���,���$�c��d��n��<mE>�9]_�,���L���fEj����?O�6��%��O&kԣ	_ߴq�%��1��r��f�#�m����jW���T�䭂��CHk��3E�ZGܸ��Z	��|R����f�Ȣ q������?m��q/�@���i
]2/�����ÔY�ެ֣&�9p-Dj<�+�}i �}Cy0UU�iD{/B��-�x��
_bnI��AE�@0��[H�&\��h�T;SV���_�x��N�����@v�X�V[�_�b�>���������z�
�s�}{ҋ����<��7���(`R�-�=|\\�/#�`Q���-�F�ٮ(\E�������<�������J����ey�Ks�k��R�l)��ֶ��!jGV���s������{�/�^27ܯ�|!��y��H+�^��FLQ��.�O������:�-�.�B̟����>����$�]%�l���/k�X�#�O�����H�a�.��8�/F���]��'���Ղ<�8i���T&6`p�X�}$��N0Q����'�[��̶Jo��q[k�z� d�	b������ L���?1��/J����QM@�W�{��s���"��H8��碀����EWOo�
_���3"�fzi���@9�s��{t��$n��U�e�1�W]4%�.�P�
ޮد�ed/���������]��8BC�����{��d���@$���f�	C<a�[��f�u8�>�Izc��$�Z�8^D��zRS�Pd�;��ڗ�x�6�L�O�o�Vz�\ǅ�i��k9�&����z]z����v��t�������������&'(�T�R!(��f�{�xJ��,nO����D6=%˩���~�ͥ�H���O�͢�唋�'��"�r
�lZ��D1~
�8����.��^�@�?���� ��M9����4E�u�{��9W![^�y-���9�F����ݙ�l�n���(5?v�����djp��_Xf�"�5R��C.�H��q�2͵�Lw)��e�d�������u�@�A\>�:�:Y@,Q�FE������T�5ފV�x|�;�S[�ɣ��>�4ku�FuwO��&����L��~K5g(<P�����梦��T�v��et�a/���'�og�3+lf����F�:]L��7iU���m��c3�R2A�:�o���Na����\����+xQhY�]�/rl�;�L��h�I��cٵe^P��qU��6�8�3�è�֐�ɔ��.�u�=of�#�����K�4��# �Zii��KVSEZ�b�2�O�҉�GQ��ku��1�N�dyq��;0��3����߮��Ј7���T�O���n.҂|]z�����U��W=�<d�����{����ē+�a����5s�O@Ȑ��3��7�Ot���ۘb�U�P8�c�.%��>ȥ@�C��n���GC���z���D�+�X͈�W��t��Yp��*o�$#�{�� �����݅8>����oQZ*Ģ��	�o��d.Jt�+����	�H.zTw��l@.��'�S~[D��v@B�K����P�ҏd��F*"d���0�ICP�Ni`g4�QHa�IC����S��~���no��$U��ۜ�_1�,	T��������^/ӘJ���A!&GRT2��t�0��u���s@��	b�W)9�[�K��k
7�%X[������Fg��/ž9����L����}C��Ԃ$�m։���<1���c����jA��=��3y;hƲ1�������G@��`xb�i9>OK�T�k ��ò7�颾�ט�'W�
9$�'6\�����1Mޖ�`7^֭���v�ʏ��F0��gt0�� ]�=W7I[:m�ɥ8A�F�nI\T"�>��W���h��Q�	Tl��a��^/Lwt�:W]j�X��ly��%}����,�I�~V1��ܫ�_@��l���%���$�Ƥ<I,S����#���ꁭk���y�O2��}R֜v��y��:i���BǌŮ���%@��s��f�����c�"��<T���/ 	�םL�ЉE��BsiZ���
���tNz���H@�%�S���������&Z��ې]�Y'���9 ��Z��^�ut�y88?�`�^}��sS�T�e�C��E1�G��@�|����|�o�[ȼ���������S%�d��VFp|�T�M
f}�6_	�yG98��L�@E�❳C�Y�{�{�'�G$����n=u��d��֞%vة��i��+��u��cPR�Aaa�V_`��pGU�Ws�t?�r���גU��f�-�-PX�a�}�*�c-r%�V��yMgS�Ӡ�c��^q�qǭq�nW�c�щ@��+�p�*rξ�v���/o��\H�x� d�((���K�׉���͆�̔��4����4ÃV"��s�Xe!������zm�qB�����&%J��}���r�р�4;�lB�3j�Q}��5��4���v�C,U��5�LD�*˛�(��6'ar��A�t����S��F�L��c�-�oz��,g���K
!�|��,�,�:;|�Pk��h����t�$l��Oe��R>T֍[�W	�������)�O�]�e����L�ds����S���H�[s��1�!Lr>/��AG�i#�Ey��%�@�2�t	$��xܦO80eΧ�Zpj6/Y�<��κ�t�A��xx#[k�\�d�)Q��̫󫴄��@^8� �r[��Ů%��\�ùz���d0&&�������ne�;���L�:1�5�]��B�������6�D_��[�A�۷$["O�nHQ�i�'ʹ�t�f�6�|�U��"��}g�F0�z��:L�M�L03���sc�OW����
R1�[�� $�~I�K��1ˑ��;��Ń�?!#;G��=���Á��	 ȯձF�ze�\��,���Ԓ<X�r�V���b���n�+%�o��Sw�2���l�ʽ��!@�<X�W8��\�EX��<{�m�~n{ �\9�a-(���� ����kٱ{[��Z�{�W���M�Ac�[��mR������S%��+�6�`�2�ӭsJ�~������Qm1����Yɺ3ҿ�"�ߒ.c0��vi��ю�*]�b�2����e�0�4�;E����#v"v���)�m��l�z-��rQw�%97R�����Ie��0�Gž��%���*G�)�~���+��@�~�`K(D�w�k\�(�H�I3��R�I�/$J�d:���~*[X�D�E�\���b�$�|ϫ�n�ɞ�i3y��I������>�O�0\���+F�&�)�v�ۼ�/�ڟ�PL&��q�{��zԼ(iP�I]m%p?��IFl��;��S�8`ߨ?	�yWK�}�2�/t�^O��X��6�e����G)���詳�>C��ȝb�3�m�t�i���� ;�U��q:@P³�1};�s�z#3��RO(19�y��Q%���������gF@c��VX�f��S ؠ�|/�� ݵ=��0���8�)�>@��h�������H�?�l5�ccp�{��v�
8{5�V4qⲰ�V�Nf������O��H��T� ,]�j��2o�����Ϥ����m�(4��-�2�FW���wÏh����&�[�7��^`I+���xgo;pX9[����XW-�#�L4��T���ڎcBǱ2܍�1	uk?�� � \��{�8�ߨ��}Иo�1��j"�R+ p��βn^���A�;ث^��<Mk���z���6�na�B��
���#����E0�xFo;HT'�3[]�U�L�V��-%/�7��^��"V�̘؍.W���5��4ͳ'6�f�u�&^TB�-���Z9�I��68o�'P�R�:+��إAxk.o�����mFT�W��">ૈX���p�K� �_{t�LB}g�zG�lL�h��U�G֖x�С���{�:ye@�H���t8���ح�vX�GA������."����b+������E�<ռ�#����~��k����zW�����$��;�j��Ϋ׻���ga�1�7pͮ��r\��d\�Bp0�3�<x�?�5~IJ��E�Wwo"��l�-"���Q�x{�N���scK��������㗘��5�4��/�T��8���F�״9K�(�_���NZ�d��H���'��9'a�$�	��:=��blҴ_@7����� ���]x��m~�h��j����,�d���~�Y��>5�u���k���<�rݜH-C��4��&_�d#�S�{�<�l����S��9u�)5 ��L"
�M����]��IC0+�^�!;��>P���aOx�H_��]�_���?��(�?�^�`��sqIi�>M����D�.u]=�5�tk���+v"※YTo)��M���4�7���I��}������-�\ar ���9��7�b��/����q��@[�_��-w�`�h�`ZH��̇��-��G%�h�`�����ڜyĥ�7��g0�C�`7� ��~�����|�f���m�Ƽ,�4sK�������QЕ� ��K��-�K�:���?%�3�6�L���!���um���]?e�#�/�wuE�7i&jm�@��_ݮH�5(v.qG-ըʰH��֥&ᖤ�W�>�w�ll�Vԧ�;�ro�⦷nd*2F��ާl2�:h�D�ׄ6���e� ����ULެ8��g/[�ݣ���]�g���X��#G�jܬ{\zR��������$-qZ��ZGXϨ���L5�U�7� x� ��C@MJ�������|��|�������6�z�Y-s�3&c��L�Ct&���<?b� ı���9?���xP!7 +/�����yN�&��W� ��	����|���&�/xZ�[Eԯ�S��N	�ifA��Y��]���Ե&��6�4�e����N��!q��`��sN�$�Q� �xS
G`o.�t���>����C�DE��ȁ>99d	�0����x �EGKe���qQ#���e�e��Բ�D���	�W�#�E��������L�������h�`G/��l���6�O[w��[�Z�F��ٞ{b<�o�Gw�/P���zK�����<[[���@ {�a���P��C��{���EŜ��k��=����bi���U��Q��v���dd���s5�_��"��$Ȼ@�~?g�$�7/$����'�8[���roI�DiR��b�?���5+((�j���E'#U*����	ƍ�iXcDR`���&NY_��=���
g��K�(��.�в�=sr��}�G�H</P++��È��1jsW�U�Ͳ������hn��L��?�������;����' ��_��b�f����]�[�0��\Bv�	0��si�<�"�nD�n)kH%�����oe�* r����Gk���B�-��:|h��#gs{�C�������e�j�7�(ŒN��G��dK��u���r�}����z������x�m ڼ5P~�O��v�����������j+53i��hX��8��Oz����a��K%�HK��
Z{�=(�F��W6Zo�$�1q1�e��IK^��w�1�m;X��-�j�/:#XiT�qԣm52]�����Z�s2��[73?Ho���`n���ijh�4<n����&^���������'�8���\���~ku�M_r��q��\缥P����~?&��M����t�[SSop,@��Z��Ab�&�3_��"�R'aݣ�����%�}Dn-��n�vk׺4&�t-Ad6a^����>g�7 �q6����;H�2���gu=պ�W�o:*�k�%A@�(��5�u��Y�9�o�xQ`�J��&�������[���*F����3��c-<�?�������/�o�Z�7�����q�B]:?�c�W3&��3������cM����*�;�����1r5}部U������: [����{F(���s]�&�vs�v ]�p���v�^��-����tA�r'r�_�{r���<��Z�&_��B�!�X1�z锂��a���]99�~;��l*;�$����!Ab&x�8��d"sK%�V��x)6�dv��>P��i@�R2�Z��4A����ճy������_�pc��t-�󍑊�e��/j 6j�����:jM����|�����(��&��AX��:|�O��sd]�҉��zhS��F0�]\�{=� /�A�(@a3�ą�0�sR�w0�7�����Q�c�҈.*5WY6o��=%�3���$� _��S#ڡ.$*�_�O^�jަkj�7�gRLF������8��#�G���J����E���Lj����g����J[��!�+?��Կ����o�>�i�[���Q��X��h��F�+��fp�Q�Q�mO�������Y�t$
��u�6�u4��mzd���d�I~��.CA�.��$ֈE�*�F���g�9�Vƍix7�d>F�[b�7i�`jh���i���k.z�W�/��+)��>x�S*��s�z8z~˭?	>��8`�FA�E~��}���0�r�?��)&���^��+�	8*9 �G$
f�Q���,F�p���!�@��]k�g�vo"sS�}d<n�q��#� �{�+Q��ݡ~��/�g᯻,}+���'�ۓj>e�5��SdRQ�G���<r##ٌ3�����7kB�
ɒ���{cK�s4�`w�G�%��g^�O������l��ݮ(�y��V��*Y��d����k�&f�2��v4����FXt!�݇����,W���7����+W́�	�O��r�EQ&�~�s5�54;�LA�=��O6����#mW=<�w�:�bD�	��J.�-�ȣ�\6iyxc
�ȋ5eq�h߯�r3	��_z�+�����אay�Jלj�E�+"Hm�8k^+��˯�	Q����{�k�	�T�G���
ɞ�&ǆ��a�y}��8[��?�P.�����}+?U!�<շ�<E.��u �2��̘̾DN�"+�W���F5$ky��0Q"�f�?�ޚ����n��N��9��N���<�e��ohz�ʅ ��l_,c{R�~�8���$��DWK�>I��(�
����)R�6T(����mg!T��L��_���L�P~��0�w�T�@F�8j|����nJ�z�;�������N���:k�驈qbBFu�c��IM�iy1��X�V]elR�f�S&Va�MH��`�2� }l�#��v\0���7����N��?i�y�����/��G�	L~�a����~=?�K1j��H���´9�l�n�!E2�}�
$QHT����nC��M��c������Z!ߗ-N\r{��������5d0%�1\��v�#挅yW�_*vοtI�g��
~��4�i(.�����]�a�ѴW�.����{9`1B�Q�pcfi��58���0�6��M`6��R?a ��vP* �d"�����k��M�� ����h��f�,�� 5��Q��&�ݣA_K����Mc����:d��r�����~G<�Gc��YZg��f���R]�*��p��%R�vs��]��n��R#1X�W�G��YS�]���:�L�G��٣yK8�]���K[D���p�YB߭�Y/���~Q�$vL w�+��w`�1���^��>��Lν�Y��-/
��!Z0n��' �3�� ���Tz%r0�ԹYH���Z�=,��=�!��{+�=�c�&��;���e������Y�� :]�]!���!+L$>y`����g���MtFCĚ�*�-��K˰S��d��i'|u��%6.-mh�����`��>UH�#m2y��Nn��kh�0��NB?.�6�Y�+���rho%(C�� ����v8ub|9=���jl�i�w=Ꝟ���: Ŭ0u�4����/�j��F�ڂ��i�Ξ1����g}0�T���\l�P��7[���cخ���%&�x)m�2a�3X��V<s_�ZZ�G슺
��r���㰳g�ʨ���c�F���R-n���ڵ6�������8�O�sNI!�>��Π7�*�gm��#�"Zb ��[�S/���� ��CgLuXC8tۜ8��ߒ��f��?;��t����+����3���e}�ܜD��H�<�i�wr�����N��yt?O�ܙ���2�A:Q|LEsȚ�=O�Ԩ ���<o� D��V�:�>}il�k*ۢ뛔��YƅM6S��G���2	���Ñk�	��)�����,7HY;� �ƑZ\&ߢ����A���m���t醅��U�g�t��� C�NP+�_�� }�3 Z���LR	����5�aRV�b@�7�ov"��-k��6����.#�0�v�r9w+>���9�"�`j`�:/awh��82��4���N�@��v��Q�n{�{Ԡ/E�H�;/��q#�4��\8t�]	d�{W���PgR�J߹��@aG��b���^nڿ�f>Q*��p��u�OU:ri���?��xb����Z�(A(�KɒM3k����?�0�97�;�F2��Q��!��,r�ǹ������u�����hX�Jn�V�-<5�����Y�e���):�8'f��fe��ls�W���F��'b`�W�����ocX�n�J�!Ħb)���liH�%�.�QA��'S����v�\IM!���:��ᓌZ���l��6�F,���z1
I��`��,�i?�I���0d�̂ol�Wm�����_L������`f?FP>��3����C��<ј�Z̨��0���.�7���X��tL�Q=����}�+�k˭=�����m{����G*2a-?�MV)��qC�e���~�S+��};�a0��Ra�Djo��L�J
2͂T�N��P"��	3f��.�TMXY���MS���ZTm�m�^T��u�dHD��o��Ԁk�w; a��[-AM,I�~v��Ŝ,�ˮ�ӟ w`�j��\v
����/���v�V=1biR�RO:�������v��lG�l��^�0Y"XA��r�Ye:U���S��"v|��Gn��KtZ��9D �ID}S�27�co+	X.!�9�����_,W>�	Sx[���a�ʹ�����YXjN׿A�^4C�Q��>u����^�1�GC?�&�����5]c<��B�� :����S#�Hk|����Β��H��T�7�/ wvя�z*p8f����K1`�d�B��	�ހ�C.�3�tǱ���:��p����8p�X�wt ���yl�����c�3hX���3C�M�4��4�� w�}�F��v�����u�	�8�9[��'�|~tun�@��1�n�Q\��4�J��	��uC�1����t�%��� ��Z��\��W���]%w���I��e�$��]h��mA)C�E%����l�ܳ�v��n&s�;��/�R��vYN4�ȝ�ve4��x��&�"���u#���25��/_N�S�>ot'ULȘ8r�O�BX��>8S�'LE�1溛�L"j?OI�c^�΀v�p]�Y#��+�T����Lp&
�~���P��=�&�:5#k!{p��&��[Z�`z��Fr���I޴[�-/��j��)Vw�S���P� �"�p|��h���O|Rr�� � 	
@���|I���i�gE=����QE�"��#Pv�S!�-���X�A�}�+�q��������El�H|s7�+^,�A+t� ^���[��1�ץ�@����w������{{O��S�SףPJk0�SP'�W�B�p �O#��j]߫&�*j�Y�����%��<Fr~RJI.%Сĸ�>�\,$��"=�?�-1��rv�Y����yI�A���k�?��%��bo�x�ĒWU�ϧy[��i��2�k��nK�S�{:�]�&?�`�����]�T��F=�2�P��{�ĸ|	���:#����t� _/)��,�]�u2�g��|�h>B��~g�C)(�A��>�g#�{K��֞�I`��|=z���]K�B�����R�va�X��B��y�<ѮU5#�N��O' �m�:���ދ�:��d�~�c9R�����پPw��,Bן�P;͕@�}��46ZjJ>��e8��s8��-�E�*���-�r���[��N�3ֺG ]c��q�s՜k*+/�!��������H醁��)���6=h����.��)� �c�<ʪ�ԤK��ty�6���*���Y��S�3q�_�wq�}p0ʍ�P��Fʨ!n�2&MN���z�TD"W�Y��s�eU}�,Ǥ焆<9�? �G4Vͥ�b�$�p�����a�B͝�۟iȖ� ����>��������؏�J̉�]ɷǇ��#:Q�:Ԃ��������O�0�;z�?�\`Z;�?cͪ�Qi�zR��[
Q&�)��)�f]5��æ�H-��A]���W�#kQ��:֌�˿�rc�q�T�]0�ߣ��
S�2<#S+�\��>.�k9�DF��Ų��V57� ��& ����w��S,�PA���z����.���%/�����I|�*7��N�.�����P�t����/S���3���[����qm�� I�c&��������20�Ǽ�*:�c�-�9I
N�-=��=����'�Wm�"?�8�́����E���,)f�)<��1��~�'�v:gdS�]��YhѤ�>��}����ԣ<�Ei�~?�kԪ=w��tg�ZT�85OF��0�IJ_�{b%�J�x}/m��[��
NH�bǭ������Jt��rՏ�;��+�S�iX�v����	k�r�j����큈K/�\�,_����y���Z5�N�|=j�q�#���Ih"��_�<��'�H["��QO��@�Ly@T+��owNd��B�2:�S��IA�%�����3J�l�'�6E�s�v3�gH���]r��|K���+\�1����]ɛ͍�G��lL��a|.���g|����Q8Vv�L^�7���I�P�o�+�oklS��h���AJߓ`�7�>�΃ۀ�V	h0� U["B��)��%���ލu�ҽ�kR+N��H���.�z����C�b�?�Jc���i�F��N�D_XU�5PؤSW�$��u*��B/g�#!�?�$���d^��WJYTN��|��U�:bN}��`<lvi�	�]Ϝ���%��E��V��GEg�m���)����>��2>9�(�;��&�U��,�����Α6���.n��H�(߾1�"_ϵ�"�<E[�4�$�D���=�;]�"�rU�I�&��d�o�䫚��B��OioZ޵������|[�Kհ����Z'Џ��:&�j<FW�������O�"� ����r��M��;�}FQ�*,�택�eN*gA�JtحQ�=�D�8Y�*��B�s���Q�/�YsL�7"+Θz����@.{���Y���'}�#��<q��o�������c����o��Cu��x<�u���螺�"�}�x���蜉�^��K�Q�14�Qb?<y���gcY�B�h��>\��x���ɸ�e�Ǽ;�JAZ����.EAMV�/��V�S6��>�,]mZ���I>��j�u���o�⳷(Kj���?���꫶���!S���v�Ԙ�#Z��B��ׇ�ؼ���I\��q~X8�ِ�(KƄ��^�,�a��7���������$����Ǒ�#C/�;�b�u�⏏	�VwK��������*������@�BZ��?��?lz��ܟ���<�Y�x�ou_?L����i�8�k5�ъ$*���zF	�dz��.>��uxF�WqS���sۻʹ�1�Ǣ�aO�� 7����C�]�Q��>Y	��F�ğ�6�Kߵ���"׬)���b��z�	��檷2�"8��l�F��e"��d$���T��I���%:S��`%6,��Z�p-n�O��� �R����l�Φ�@? �U��3t"��P����R�@����\��.w{�EJK���=�x5u��Ͽt��S���+�@r�س�6���u���6����1U�X�����l�o�
���l.C���'M����{	��ǫ��;�A�XH� �*�h,k���Z��$�����v]����3;@o���xH��ya8_�>ىY�'��"��[3��UΚ糼�E�p"0�YCt��h㳣r@^��ݤ�<A1�l�S���&F*�/�;�N<8�
�W$��B�:�崁,^��;[�t�皐�[+�:��6,�a� lM��^[Z��]���G���#���L&����������;`T���8& ��7QrY��'{`4�Z�_ST�_ H�m��o#�wFe�����}"������sP�u󪊀1�4�cu�2>d���nnc��(��Y��+Jo��}I�:��gX�pP�U�g&8��=_oLdr�%���87�V�ZC[���y�^ˎ9Ahk��Ny<��w������P VL�m���/�j�T��IC�����keQ����K��T��x�jC.Ip����BuS%�DP��b�j#��6'M�*o�*gx�bә��e<ZnYɬ��3�g꺙�Q�ϡ��9� ���݁�ɹ'��<mO���awkI�ł������<�E4���Xx;NtB(:�/��	0B�DX4���̲r%1>%x~�9u��W�� 0ā6����Āp,�Q[���7z����٣�*�i_��5����*)�}B��*�&?�Ѻn�j����^a�r^�쟬�+��5y�s�NL5њ�R͊�H�h�P�V9 ����ْ@�����o5�2��l�,��9G��!���Z�/i�2�[�����k�'��Re�3����* �+vs�3��`�azf]�3(]&��%��j�`SB>!�8XPmx�����i������ƽ5��ڋ`x�kv�+a��Ep�sh �(����jC}�f${_���P�����%G"�]�b��[M�#���2C�%Z�A�Z<G�y<7�'&_2E��f�-��(�2 ���@�/��'��<P�6/W�����:���Vy����4�y��&���h��%@�wQ�O�ZI$|7�_3ͨ�+����Ɯt���Ur�%J�A�P֣�zFZ]z���}�e6�C
��0Rlc��(���9�m	�ikZ�c�S����	`\�M����l�i�V�J�"ʜ�T(2a绂9Q3�o����>�֦��_���84�J�]��
!\�I����l½�(7@������x�� ��~����5��Z�����6-�·�C��'���!�i+���&�[,Hi�����s|���%�nB���r���58�&��L;.<�.ə�1%G�X��U�@�
�N<�{,�&��OY½!:�rI,��m�_�>�w�0�m�er@���{G`D#�1X��A��x�m0!�t���$� ~:@�
���((��i (M��?	�p���f�����?p�
�]�������1����.V*��>��#[]?o	���)��=q�*���: �Y�o��1ő�MH�;N�?��X���їr��stÂ��-ܺ��)�Q���\��r��7{��Wu|��:����Pl��/ډkT5+ֱ���܇Дa�B�1u��0��gD�q�T�[��
�I��A@&NA8�a�o��f����Z��楊��k��⇪��G�j6�䘠y84��d]3�]��R)g���6�vA��r'��8�#9ُ�q�=���׹���F��<��8����c>�;��0F��3�5fywMy7�=��kQ�>�g*	,[#�~C�C��P�I^?�\.K�أ�Nv�@�7��-�Z�}_�5��T�,����`�@(��A�4Kx����KzI�k����q���yŁ�*uc����8��t��ߚS2�a���O�+��[�&�7o I�M����d�G=�q	nM#�a�LJT󒕭T!6q�lf�� 6���vu<��<P��s`V����bNy �,��n��5�&��4��R:�9��ZkE���>�w�ЁB4Ų���Y��~��L�B�������8j	��Q�������(�����$�Q��%A��P���mCƵ���5S۴�u�2O%cE�=�R��3��^�5mˠK�|��p�R�TgY���9��yPk�:��r|C�`-Tw{�u�()`m���ͦ ��+`77l��k�h����$�5���ܡ��&~�MϷP?�pݛ\z����0�e��1�)-���#;F�o�{�����
�����!�fj�����>�K��2Sr���!�(�g���7i�X�畤:���������u�+8���˶���*���a���?֥c;�wIf[}J[����A
������ ԢYs�uH�]�/�Ĝ\�f%�9�I	���)f�žn�it+4J��+s3}ۧ���l���F�� �Z�Zy}\{�|ҝ�I�=�d���BU�@��L8L�񉯶�!F�����uR�ոq��ٞ�����@�*W��E�z�N[�i�{~=���"er�7AQ�>�?�F �֯r���%+R�I5�o[u��f�8���DY6�29��rе9�K�D48��✲���Ձ{�-��MYh��Z��&EbØ�΍@4mP�э̷8���!5aK56~P���}�w���'?�_�3b�D�A�^=/j���%D��|��v���K��*ЎP(�n��4F�4��!�(�ש���w��n#�L�WN�.�Ȭ�\Bs�q⁼= i���b}���|/v�T/�]x�Lz%U��iT���xlJ��In��0�HIM���'<�͓�����F("�F�Dِah����1(���	.vs�&`��t ��G�m[�#��'�����=�Q�z�a�/߉;��K�~X����-��z[�V���k�4����k�׎k�h\��&��ܩ�=!�V�_�T�u��N�S;�3so��)ĳ�P�Bz�rTi��Yp�ƀ�/�s����zu|��Y�/^|t����3='6�NH�fJY��2@��Rv4���k� I?c<K�2C0���˻�X"�A<?�Dܪ���kZݻZ�P7�%�2/����'��R�6KjE�j��� ,�C���Zau$���$��qמ[��W �N�e�_d	dƢ�8��a��x��e�X���h��AA��4ׯ� �1N ��A�a�t ���x�ک� 6�{����;T��-�_P=�x�-����Z�#a��'�>!�/	Yi�á3�5S\���6��|Q�&�Ō�˰��h�9�]�V�8E8SXeCEx�*G����j!��&����u�\�)7�մJ�&�D\�wn�Ո�7_ema�e���j�u�D��J#��l�L���*&�x
�1�:��N�1�]�5�� �
rq�u�o�\$�|o{�G�
"'���P�[���c�,U���ܤu��		3��EY�<C�@��o�|37N>n��((Tw��}�*%T��*�M���7�|������I�{!-�;�p�0�KX�(�wZ�\������)�H�N~���	���!�s����:#nG#տ7֙��.�=:4�������$�]3̕�6�R�vu���p�!L�{�{^i�f�����Q�&�/R�ǬO(L�c������l׻'9c�P�y�I|.8����d��sA9����jfR<k�]�76HR'9��hr� vk~�q�D����T_��0�x�2/��Ix{���H��A�A�I�f�0�c�ƸA�<�{ ���?�0b�M�19����;�*b�:�7E�N�����~�|7ąNU_��U��+|ll*�"��,��~<�a'm���kzN��3C�Ϡ{�OI)>H�P �EV2�5˟�l���b�b�Y���U=���(����65�CaBڛ<3�+�wP��gr�0K=V�le:����B���v��q�0���P�<�{���/���w�S����5����
���h��D�i,�E0h5R #��5�K�X6 K �c�7�`ͽ��ȅL�J���n>T��>&���L�N��F�-.�V �J���=J�5�R��q����wP�uZC��j�놽���3�T��!G�EBCX����kZ���0:f�Wj���ڃ�u�9�����Z�F���)���o�G��T-����v\OFy�:O��e�cg����n]c}�g�u�}$�M��և�+�����F�n�#�
6��p��אA{T^ww�Ҁ�4c�G�7�'��z^F
j��1x`��l�r���$d��K�Y�]`��|��*[��%_�>ӄ�ߧ����V�E�~Rc%�Ӯ뺺ԅЯ)_�C�r���$�U�x4�+^������YbEg�I-�.�ý�u̓�4v:�n��Ԡ<�vH�)�,�jD5g
����%���ȣ�({e�b���[��5�{�j}Ѕ�@����Z��Ȧ���Y� �
=����������~U�$����^ǶZn�$��������BX���K<�,�t�4�,�"D���E?��D��|2��y����u�̾�t(�}����,�495ܝ�hd�7���~\�7=� ����1��J�$(@�,�DOO�HLV�����.]��"�N�U7��'��������	���h�z��(�@���  t8�p&�A"Ι��}�����W]Dͩ������8L�G�+Z
�d��ǥV����\�HtH �l�W�!dICA�[�P\<M%/�z���;�q�E����eM`l���oy�����A������t��~��y��JLe|9��r���h�k�e^�Qv��B��]�TӸzF�W�(q�T��%J���b��b��S>E�l��4�{Kh�i�`�PMF�+�ތ���cj7�63��&3B������r�9D ²������m�P���i=����w_)�F��)/�ﶖ4��׭��٬A�4oYz)B�û�O�;�����Ò�� _���b�f������L��ZK�!Dw�E�T�Q���X���Т��'��r��GH�t�zgK�Z�����>�0&Ci�Ɨs�e�c�9jB��A1vU������B�!�G�J�E9đ��[z��V��a���s���i(&���#���Z2�&���Y�� �Nx.�p����t4)a~��Q% :Rp��;A�\�ʀ��U�srٸf �=��=�Z ���QoMI�@1���ҭ@$(�l�l�;i��Xj~]H��Ƣ��@)��yy�v���45�����G�m�\>�&���g��3jCEE�j�lĮw0��3� ���4Pv?��Qv�ڎK��`�[���b����g�)z��".���S�`��	ה�p�!)��Q��=o��* E]��H����K��;,��+�U`��!7K>Kz"��y�����\:�s��iv��f����P���+EZ#��c7Ǚ�17d�fj޼I&��qt��L����[��Pm��e�Ǜ��.6B{��,H� \<M�>Ś��9��t�	�w���>� �S���<G�~j���E�Q߰��6uNR,ˇ���D��!&�\�h�R���-}a+4�.��]/����X����G�I �5��ق3��iD{�K�3�8��C�$��V��2�1�e��&��Ui[��&,��q߅2��1��d�sĳG0�	��&<��p��~d7c.�O
� \�|�k�S�����l#O>�l`����L�#�⁭6��@iR$����c�z�v\&?�q�drS�d���$��t.���p|�;m�jz���bk�I��W�#�������)�B��Ƥ(�H�IDw3V������V~B7�Qp�,����5����|/7���f��j����h��xǪ飆�9y�.z��)Owڇ�������t4�n���e�~��^��Ul�f��=���c�m�P)W+	�ӹ�vK�mɹF���e��Sʹ�7� �bp�m۫Cv�m��"�E?��ﹺ2�����R2z�m3F��j��guk��7ji�W�V�z,�ϊL���X�� @ QO����<��!�IFJ2\�y#��A`f",oxUb`���1&�!��3����aK���`���dL�U�.0��=�3a=Ϙ��)���>��NPcԐb�.[�� bõ/'�1�& ���񍂩�E)��+�G�N�Mj�t���x*�;���4�5`?�k[K|�Mp�����-X�[`�x�|���>�j=�~���R��)Ѥ�I2Y��pҳ���O�γ��p�P�	n\<�8�-Cϻ�)~#r�sC��@L�C����r#Mr�|.S�h'�ʌiCK�� �ƙf���]z��W�U	�d���j���N�}l��!6�ǹ���x�\��h^Z,V�c�:��T��<���Z#�=� ���B�Om��%0��a
 �QS�?^�ĵ�����ڄ����/���Lݼ<�!�ǈ`��U��jP��?�ێ�z�oCœ`U�61��K(x4��Wd0���o
?��XI(���|��1�h1�+\�� �X���ϨN"�I&����ӟ���[w14�6��E������/�EP��e�cK�`Uh��[���{X�;�f)��:��~_U	�<r[ �����!��܅_�x₝�]X_j�j�A��O��cW�����`�h��� _���R�ߌ`�l}51u{U���a��*�i���'��"|p!b_	}�7F���#ť\\L�ЙN q��
�}�|`�4MTѱ=�!�.)yI#\�Q�&+A�:�9�%�5>O6o�):8��~
�O��$�W�i��w�2����|�&�?
�skc���L�%�?��W�r3Q0/��8\���?�G'�:�Մ*B�	W��^`pz�-<w7¾\��E2x$�b���_�'�_Of;f1iHD�b��@�(�H�F���yǴ/�@_Ƭ�b���>N�1���������i:O����W�Hx�s��"�q��`d]�®�=����)����������
!��#�~8�f�د�JD��~g�� �%b5�P?��4�Li�<���W(�M�2L�Z��(�a 0���i��I���mvG=R'��iL�%2�1&��%�=%��=��*C���R%Z
�ZФ�_�|�*z��@��u���D���|ڙ�D�]����_p�x?O��_�tp@�v�$ҋX�+:F�<L���r-��:��t˼j�T�'����8��6'}������m�B�$$����#�{?���֝���Mz$��h�ܶ�Q]!JB��[��
Ϧ�r˙Kp�T �q���"���b�1G�i� 
��ʀ���d6�f�ss���ϰW�a��?�@�-u������j�2X&!�ͪj����K����b��/rx�Y�J,�y�)j�Ť���z�:�dn�dm`�#�����J|����"'+:�)~�h��}\G�V�^:,���)��T����ɠ�M��Ï�䵯5�}��n��~�Tņ�Gtߙ�}~��Qc/�]�AXkm'~Մ�L{ߙ�W�k.X�u�z~ǀ�FՐ��j��EXRr&-�[�"͆��מ2y�v�r��ֽS����S�jH؄%1W�޸(-(6�({e��H���u��Z?X5�y�K����eQw`�;|HG�%��`�Y�GpG�&w9��Φ{��l�Bj��*�FiM��Uf�6�8��~"�� !L!�Z�˨L���k�v�+�@.`��W��WJ��/�b��D��V]:���S0��,���LҤA��k�N�[=���V�"�n�+�D��c���giQ�O#���`e���U�X��@�� ���S]j�Z6L\���+l�u�H�g�Wl~�o��o*��7)X�K����a�d[l�;)Ӑ���+7��C��<�@9�R��<�ټ։�5�5n룶���L��i�Б��I
�o��M�  �Jq����R}�*����|ĤkW�Th��6�+e�9ҳ��xƃ<�R�<Tz�Q�E�7lD�?��l�OJ�:�����K��o|I�5ė�[ɡK=)��ϊ4��>�� `r��溨�j���*�=�Tꌗ}�k=��wq�˜�(u5�'�'�.�>��b��RP����$ٜ�iD��'���%Ι�[�L��Z��JAI�I�4L5�X^�`�}��2����������2ge��=��M�<��ُ���m�jR�̪h�+�W�����k����;4�g;Kf��B,�KW	�n�-�F+o����Z^����q�G
+fn}�����G	�y������ط��ML$��Q���`�9��T��9C)P�K���aUx,b�!в�}N49^ޑ����z����h��p��� ���/��>n�c�?���@@�'�z���&�]�ê�F��hC�A�|�y�;*�z��������4��T:�\��@�a�b����H�'w���D��̈���4�6X�g��OE�Z^:��2��H(����ޮ_���08ТP���N�(��u.��2�}�eg��2��ޱ%Ş��+Q��(�a��+H����)U|�\���5]V�v�,\t��s]�4+V3"w���6`������n�Jd[eo�y���<鏰3(��êO�:�(ɶ<'d�Q�#����͠{8%Lfwa���IZ:Ă�d{��J��s��F�N���_�>�2��"�7��:��K���E(h���(ȟ�@p5W��u���g3-����/�om<�,e.���AL�:~B��X�֥,D�6�$h�+�nk!s��H�ݐ��!����rZf~��J�Tږw�*���gW�6�S�+�_Sir������<Q<�e �P���CV�UX0��j�� ث�>����S�A�u������M�&�ʰi�g�(�,��9�0-H��cԜM�ݖ�
�`��e<��/����Ҝ����S�2t2Ս�����`drf�n*Z+�?��+T#R8?����,�FִE��h�z�(�j\rlX r�R����N�I:�,Ϗ�:r�9�d�@���jϰ�#�&p̽߂)J�c��G�V��2n`9����b�
<�
���1�JSe;f�	�Z�W����䂴���w�W3a�N��p�ҩ�#�)G�a�I{A s��R��	�V��P�O���Rm�γ���Z�Vӱ֦]�{nB���)�ϗm��y�����e��3�oW�p��(��������d�ܐ�7���u*-��+1|S���$Ri�w[V�~""�|v
eh�X�+e:��v"�RW���s�N�r�*m�K@��w�y���D���/ɍǚ��7&�Ɣ����\E�=�r�����{��s_��l&4�XF.F��:B��Je5�.T�T�c�R�����=̨'�o���HE5�7-�d,��#S��������2���ղC�~mS7��/�����&�E��?l��}X�8C����_R����s[pϑ�5,D6p�*<��?�OΕ~��h"���kސ�������������nvh�g����f�\c}bbt�,u=����������Q�Za`ƀ�����	O�w=ѯ���;1ѻU��Dxt�P��%J��C��ˣ�`��e�ijQ|����i,�֚�FC�f)|V�PT�/i�j��(fzx[!��� �1k~��1�p���a,���_�N�T�J�)(�k�/�)@0�({�O��k\D�݅��۰���T4h�eqW$����/aU���
H�~xQ��AtJyAL���!�PhL+�]>b者�t�f���w�U����2��n�ΰ������DKJ$����>l��u�XR}�k���& �w\���b�;�-J�$O�d�uܻ��!`�r���b���tG�<��7O��.�z���N����o-Էv��՘!�/8�P��Ӥ�p$l�y���v����]oFiF.����Jm��@�25��@�n��uM�W�` yz>&��{6^W��IF����'�#W>�1gB��z2�Ѹ㮺#��`�&}d��W'�2K��H�ͪ#�C�a�\B�mnN�4�q[סl�9����a�V�p����a�v7��!��M�dk�PFk�Gs/�|tY�g�yQ|Zݰ$g�0�Sf{˾��r!=<�7��.�ʔ��rNa
��eB��x�c�#�ݬ)`Bg	(B<(�\���Ƨ�E!N�DAE�`��1�j�hL��t!J���H�98��"fq�Q�x����l�o��p�ɮҶ�Ybq�z5�Kр�V��_�Ծ~��d	]����!�'�g�X�lIlە��y��h�=~���O�H��iO�\M_[�@1f��QS��a��
Z?��e<��v�"�'��d�Ar�A�����4�zY���Za$�>6u$F�����@z�]��FX1��=�������VZh�#��)�p���� �������o��Bu��ǖ
�=	��.%��m��IN�uI�}�sC�xQcx
��9��i���J��)�%|���7o������+�5i@S���jU��ц��an���������n����H��n8ߨ�zc'�eB��MY�!�g�"	��?��������w�3T�}��𳐒��Ď�zu�)�k� �J�Uy�2��
"Gl��X�ր����G1)*�����)�Ҍ�u���HѺ`��y��>!=I9c�,n��%��U$�@6��r�Ȇg���h\~�7�]��f���aj̻E���g���0#1�k�tux��0D}+P<�dQ�i_��8]�'j��g� �����D�4�i�ڥ"���������<�G��H2RTYTO!6C��^�DΚ�f:;��L����W���N�=`@�*d[���@�9��XR�r�s����8x�L;o��3��?:mbY�"'+\��·����\��ǕKͶs0�������ڦ�n�?���*kx>��#:b�#�b�+v �P!?L���+�Vb�q;�љ�v���/�\�KW�mR�0�llYF~�|�/ve+�ú6�9�״G4��ʥ4w������0�c�5�2��o'9�zw��\){�W`#(ZӬ变��ᔇ�0\�uW���
>gV�]�7���2u�%�ۅ���:�D���"�R������c�|�[�ل�"����/Q�㒍�J{�����.`�����,�W;�啸3��܀]N�w7����|�2]�D!/ �9�m3'�D�{�F�<�lr[c^�T=�F@� Ű���0�v��:k�Z �R��a�9A�+���,aC&���c�U���7�7N�6�`�/mؿN�¤}O��6m�((�'K}�1D���! Y_&ae�����}]����w�.v���,�S��h���3�C�^���e�K�t�}>j�ZD�{I`m�VO�����~�U�iUWċ�W�����aH�6�0K��h5t�SJ(lȝv�S�P���vm��\q��	؃n'[�5)������S�lԓ�k��J���Z���m���J�vwW��^�G4Ùw�����?�e�G1��Cw�-cH�xjX3��Ôg^n�rE�"c���z"%�[���@�Ԭ��.ӯ�QQd�,7������[�L�B�q��>~
����sa$rF�`���B�
�vr�V��]U<���m�`Dx�>A`"u�=��9¶�e��9ړ�B���4�_�ZE�����p���>�8/�Y�B�e��Pj�Z���c1�1f�)�O��M���tt fR�L*�`yZ)��[������9��qx�H��i:m��������Q��t�!Fjz�n4�c���TC����*�B,"	2�o�]�}A;���E�Rj;v����e�nW=�-7Y����b�5����qb!��u�'>+SU�>v���烕׵�*;\5��Ȇ�p���U���J,���F����HR��e�>́�l8��r�v�|`�a��WHCс�����%|��\��k�4q*\p���7��{���q��(�?)ᩀ���^�=r�����RD�c~xT_��AZg����+4I1�,c��h.��%��D�(��ag�*P�����K�b���Q�+8uԟ��c#s�W���"N��w�&�꼨OӋ,����YL��	-�E$w�����苷�&�� O=�.�c�:��"��]��a�)��x�l�"^ԙ��&�d2�nXn��Ey.�!�v<5Dp��J���m*p�56�����g�e������X݊ό�e!����`dV=�h?�wR�4X�;�E]}�_����v�p@�Z��t������ �������&�u�M����N4.�ˈs� ˟23˄o���E�*����>�O�/�1���2�C���S�M��K*�����#��QLr�
B,K�뿀��R����`��y ޳^F*��p��jI���,̬8(�5���.�&WM�T�[��'�t��A.��SN�!-�3p]P0A�j���_T�<��l{�ɀ��,����D}1���<5��=�|�B��7�I&$�_F,4��1���^����7J*4��T��˒�k�Q��ϵ**�Ɠ�!H�����O"0W��XẐv�ڜ@3s�oC��H]��Κ��{�<�J��]Lk2;p��`�����	C6Et<�:�#�����=��`f�L��(��eދ"�1�	lp���9��1�*�{,8��������<J��3EIP��6��A���&ܞ����"vp[|S����tG?pYJR�w�5P���G���(�͇7$)�<��MH��޹��h��(ڎFd!"��.p�F3�+�*YS����~�5=��j��p!g!���	,�'Z�e$X�M�-���c!�����ȫ�Y�;�e���N\�p��E,�lyA.��Uh��mnЯ�E�?kD�m�E,:����2�\%�N޸��c �2a��o�V���B�+��2���z��d@|l@J��MV}�E�'NԨ�ƀ�y��AH<�+pR.Ȉ����O# �R p��YP�ٟCD3��qJ8 sJq�AH�lrI� gf�>+�����J�cˑ�o5���"A�� v����y��:n�Ĕ����Oy�壬�ܣ�X7P�'�`�S�Q!ױ��wh����x�^��y�a���+Qk�oC���a>2kb���c^��l�eKҟ��O��7�E�M��HI�dw��������uV�+v���8��D��a���ߟ�z3���tn/�=��eecN��K��9.���4Ei��H�&����,�/;��7�|K:6�bJu��������v*Zn���(������,y��TB�Z#sm���ʹ�;��I�$��'��U03��d�XWy��<��Xgr`�A�SN��p���-)cd[l,�.e�dn�ʦ�^M��~I�{?�v��_紶h�����|���{���dd��鏗���.u�YL�/3��seU%���č��P +>Ml^�xJ#��1KV�c'
�QO3���Щ����p�t x��r�Lݬ:�u^<ql
��k{l*q��^Jt(b9g��?9�?���+�����:/,F��<\���%��V�f��$h�9��t��o�6d�,?+GD&
�9���7Įv��QKUi�KӁ���~\�"�
�v�s-i:C#7�Z�2�]�(`��X!��1ğ�A�|�	P3���;E\ߠ5�a	>�cAW]o� �.�IuD�d�	�c�_b����"�{�x�4Ԟ��F�oD�RG�`����'���^l>HwL����M��G&|����)i�+p��+= Z��-��ze"�VK=pY��f8�<XQ��U�y�ݟѫ��~���͑@��_5����Zk\3ak���e)�J���=�^�v<'���5�����5|�wL }�߄��Dl�.4��ە�o�NU�S䐴���L%y���˖O��mиDJf���N�R2/z�_N�W}�!%^�#a�~R�;��H*%0���a�F�GKh�龿e!�����9T/H�5y�t���7���15^I(��Ԡ�.��L��נ���F>�nS���]�-c>d`>Z�~�Јka���V[�'�n.�.(�k9��*�$Ο$�T�ʔ�&��5�VT�෋�rI2���Ӌ%�E������M�vc��p��@��-����0�Y��U���3G��>i˂T8�s�s�d�Om��7����Z��mTv��d�!sԋj	4�d����g/`q)wB0�;L:�?ˬ ��Ca�i]��X�w����t-,�S�.P?��v��7PՖӏ9��nL���3?Vw�7q���?� �!�%�i=(��ì�C+��ݕ˒0�̮��m���/l:��E.{���Khzz^ǙI�R��.�k�ץ���"-�C�%�u:;[�ɛ�JH���o�19;?� 6!�7����z�,a�{�yv���Ǻj�	�9r�k�/`�D�r��:#��v~ ���r ��n�&�;E�S���͵_����R8]>���P�|PG�}��tPC8��Y��Eg�m͜} �h��yqy�nE Lb�@'Ue?��l��sd>&�:O���o|��(��%��Ў�H�*e��g�_@	�����<��y��sw�k�6��?B�'����R"Aȱ́�_Bu+���Ti
�g���s����C�V��ߵ�]�����K�A�I���Β��]01��Y�Fb�B� �	j㐣zz��U&�����r҇g�������9P�<���?��iY&*=;�����}n��ξs����MZ��~��e�vr%�~�1'���~G�X�(Q���׈�/4�q }�i��k�wx44�H}��-�!5���
���5,�y�[�Ec��Yo��c\4
u����]^(K� �A�@H��&�t�3ࠠC�]�|E�ѣ�7��S��J;Z!���"?bC��`H�� �~�hq����;�4���΢&�N�쩙X��A�bؠe��OVJ�Q�,oy���d��������7�����;����M1<e��q)���p��%�p�R!۽f�kT/�@a��-6� ��_�Z��wٿ�6���u#'W�NyO2W3#1��ДØ������?St#�d��n˟��~on[²�є}fϵ��c��.y'�����n|$\R��j�����^�!�0v��=y��-�ϧ�q�]d�H׃�)��u�co���
��F]�q�M39M��<:���]�8M�(f�N�u��ض%ب��M;mm��ǽ��\Qn�򩞪��>�����")<�@��Y��@��Dr�D W�����I�R��=��0����h��6�0���f�]�f����ּ�2���Tl`>7��%�8�[_!�^�s+�X�LAۤ�6F��w��]�y��YnZ�`u2��G�Ωg�&��ϗK'!�x�m��&���q�9\A�clK7I��ٲ��j|P��U�p��3X b	T[�k��_:t���Auk��F'H�S S}6�Q��AlA�3@��@V���3�=R̉A_��;�;!n'���w�)h�x�se5(���[�ô�Z2�JU�q�F��(��!{�X�K�H�7	%v���0���� /j��xcJ�y[:�!�dE�[��1��-R�>	OV+�`��O�V��S�������cV�2�a�S��k����!�qƦ��ʰ �O��b�İ�`���ԧ̢+�2o��i�!F�)G̪��/׈�9���[�׶@z�R�q-�t�N5��x��i�D�.�U,Y�<���|���-�ªM��+l&.�Sx�%�¾�C���(����?};�3Ul�*����U@��+�Eǘ7��E�ݬ�δ��%�Dq 2P����)��io��r�1PN���a��#d�M-��";�`c,7q���	��bS�!�1������3|(4k�$����=���歑@�"�n�2}h��G^�*�U%��B1��=4i�xɃ��ipAd�3���~$ׁ߂��GIi��\-��t���1��F&Lf�'FaiB�"�]7�͛���ׯEx�E�,���J����~TV�/��X�]ַ|��2����Aw E�m���[a�c?4p(�,h�+z���-�������h�Eu�_�$ aS0˕�v�p^�u�B;���	�sɠ�����(�3!�uAN�m�(����8F�luG�}�NN��[xŋRo'�Rr��hy#-��ZgyE�u���AY��G�>I~���@�`)�i��n�Rb��v��x9m�I�S��#^ꥉY���k�Km�ш!�T�!5K0K5K �ל}Oz�3���ɔv���m���^��:;㢒�]�y�N5�]aqϙ�5X�5�6m��IX��Dô�j��)`"�gH��//���֗2c���/)������y�W�[��V�����Y+ع���*	S���Ukr�y���Nl��,w��_v����V��2"hv�Y��T��ؽ��U���D��C��7���2��۷�����p'�Q��5�i�L�������<В�����C��fш�Q��{�b����GzB[N�&��,·�C���B�k��0���]}�5���b�9%9S���g+�Pnf���lo�5S�(��Ӏ��J����\�h��\:���$0+�	�/Õp�@s��:G�50��]k�~���=�}��RR�C�������GOf8�YL�![��-�҄��2����ڕ�19�13�6S�[UBlX�ųr��g�s����ƵVK.sDwW��d�$\[�0�f��W	��"�;_�jU��� ��7.�ˣ;X����d�*��c#�mH��et��?������hJ���{ݑ�AG,SZ�L��j���\M�5��q�q�z�[[1z��S��5T�i�U��X�K)qJ��m�� �-�}LE��Z����q(9��hK��U�s@0"�� JI~��DN�C��<�pm��Ǹk�F�PM��(<��JB�[W۾�J�ц[��!o��ek�+�u'�w& �$a�=`�N�l�*x�~<k�ل+!DD�x]�IN�렕�2����1���qx�%�u��mn2��E��:\ި��C���f�.V'��Yh�'��mB��Ry�Wg7�H��Zz��ۇ�y��
���1躘�l�;��'Z�)�������C��]c��`Y#XѤ��RP/|l�����2J~#{�ka��dۼ5�,���9���O��VEP
�9�
8�c����ղ̣�5��W�kY��9���!�����*��v�|l�#��D�c�����̲�w�xo/I�LfLF2�h婌
J��l�������G�X�[�@C��Ύ�x���5b V����	���/\Ԫ+��M\�l����Z�H(R����)R�H^�,�%{<�L���(���M��r��xR5���V��NCg�'M'�����1`��N|�|	�r��������js��Aw���g�����iz�}7�� ��{�{����܀ �u�"���؞o�[:��W��ʘZBl;��"�wiL�y�Kkd��wa�/.0�y#_��)���+}`�!�	�$7l���f��䏺Ҁ����X�"ǉTH��XC$ޭ�+2qI�ى��먹�a����|��LT�B ����!G�-����/1�6�~4�Y���C/�Ձdt��^p�Kg���.�X��z�k��"`0�43L�a���*�[ku�ɤ�U/�=Jg�X��l�ϥ-Ѐ��W�j%۫�����'@�_$�7m��9�{"�"��Lmp5`~_�f���N!av*���o_���p��E�5�ۆ�qϳg[T�G���݇u��(�g2����$�X���k��얹#-|k�4 dЖ���_�E�<�Q�tR�i���d?X2%����ZF�}�m�'����(?��:����\��"}���U\����7�S�DC7Ӆ��w9z�L�ƕ�M�*��X�A�A�N��[u��#X��O�¯,V�G�e�=b����*Hj%2`��Ϋ���Y��)��yF����㭛��.�M6,XJ[�{4qr޺ ?�@�CP��zTI�Q�}�������>$-�z�~GU9��YL*���ztP��B:�s��s�+�A#>����VXA(����;�������a�+;T<ʿ�w�)YQ@�؉ �G����Ds+z/���%:mv�@��(��Pàma2d�F73w,��9L#��RL f�q^�5aMx�4o<=dm����1o�����I"�j��D�s45��0&�7�OP�ű�+�R'3U��`�u!O+����P݌?ai�Z��x�[���]���8!6X���]���bu��h&:B<DՔ�8P�JN�r#"Dq|��T�V�� �"p��~o�!C��B�G�8@F���7}j��)�e�gI�M�=S�G6NJ!�j��������K���;\��>�t1�2\y�h�a.�T+81���(��Au1t�ɴ�з��}Z$ƣT�$����=-���]��^~����/L~���g����ˌW�suؗU�M�o��4q���A�����q�O֜�R�B0���.��9>��[��t�ml��]��7�h��9&SH�Eos�v�oi\���K�D��}�D��N뷳�L*��R2�(�_��@�q�q����F�j�P �FYuJ��7B� ���ۈ�%ޙ������s�X��rA�Y`���}���K���I����#�ݫ�7$*��Iܟ��!E[����-wob�f������&hY�[Ce]Gj'���꽮W��8����7�\�J����&�ކ>;�ܞL�T&��%��(T��ݣ�o��P�����t�8����Üf��9�M�@�W�a��@���67��LOa�:?�I�3��=X�u����~���G��JNG�t5xܴ�@�'B���ȴZ`cO�s����S>٧�W�y�m�$�����͡L�밆��@WicSs�"�^pM���
Ò��yZ�b�`�<��5gب�����T�W��vW��N��$�/	qȊ�@w�%��-�k��p���w~[OS�L����<d�a�z=A�Ҷ�J@�rW�
�Z��q�yLv�1���
V.�ϧ���Z��g�)�ȜМ���i\�۸I�9�5P ^����`О���oy�h(4c��kE���"�M�j��8�;�)���e	T@�I~y���Ȩ��0�V�B�!�;���A9�4a���_��h>�A�����OǮ�3
�[�n�x!{șO�Ʒ��kj�#r�����g�WF�Ҟ������K338*nh8�ܿ����_L�01=(��	G�f��my�7��Ug���$��$�� Y`��5��,��$�	��"���!Tƿ�(�"������G�q����`��c�~	�r���;{y𱦓.�%I5i��)�e�X����I��7b����O@��bZ#Y=t#@�	�D��_w߲�����.��YM�5��OҴa(�zAn_?�jYS�(�a.@�.Yܚ&������cpG4�JA������9}�D�Z?��V1<�t����+�<gRl����������!���wոy$�x��@F���,��I�]��'�O4�l��rMi������/RZ���Yph�!\��̱�B]V�P��w�ů��B��z�ln���G0��*[*;ۙ9NΣ���ڷ��9�F��g:�i�6ѽ�1��/�w������hs���g����6��*�����<����S�'���H���O��~��̞Y�qpy�ݘ$
E�7�������A���ړψ�&G��f|��ov`~��$�7�������B��S�/���n'_�@�q�#7Έ��X��?�Qs��+���A3d��Cr9r9,���W�t!��c��K�>��AD	|�2�3�wI�_U�~�:?r�C�`^�<T.0�;���̏ߩ��X�p�!s�ox�y����ys4�ތP����a���<C��侑qE0n?m�B�X��Wl�����XJf�
2�(�2��
AT���D����g�p�ՆZP�k��f��0)oS�Ŏtq!ћe�j�k~�GB!˱���ب]\2Y���B����P�WQh� ~vH��H����Ȃ��.��mxN�8d7g��2�gGk.cMr��רF2�&�_ON�2-�t��|m��<��3�exQ�/:i}�I�.�ՐF�%i��d��`?-�A�*!'p�v�N�J^����WNz��cR�/[|�z�:Yn}��;����NIú2HV��=ZץSq\=fP�\ɟ ���3#�<�ŀQ?�F�]��;j�CQ"��K?ܘ(/��+���l�����b�{���O���G'����8�w��}���7��pz{�.�!�kR���$$(���)yEh w�����z�\^��S$�Ev	�U�{c{0N��[�Յ�7ʸc�;K���1S�'s���V�%+�M�tn�?�6�2���ے��f���,֝%@$������~u�����q���`r��8���em��U�����oV3�Y�)��;�e�61�x{S@bk�f,�y܈7y�6���%�-YIO����of������ׂ��7bX�S��0H��NYK0c������M��-vLoC��܈X���1�1*�%j9�����Ь
}�{L�����-�V����C�� 
*Y�N�_�C�D�ap�b=�[i;���:����b�!�~!U-�Y|�&��bFG-���q0��Q�.n�2	��z@u{�Q��F�fF��F��t��Ml+:0�&Ӻb(���Eg��g�lbu8��U"�r��S��q�23T�ϕEՂ������tQT*�������އ�hO8�S���]�c�r>�.VQ��~��1�g�Y���r�[�T������$?������3�H��6�k|������������|<&އ�z��m�vş��Pv���[�u]`�ˣڇhp�ۄ�g���'�~X��Ҙ;=*VMp���s�<Y� t�g��*��#����0�G�I��ֵ�Jx�4!��zRz���g0�zt����S�T������s��>L�Qm.��b�N���y�Eۣ��lM�&�#=!�b`w��q?��{���z�OH#N��l?�k�J�T��0��Dzz�8܅1���^SH��(�BR˱8n�q?�v�؊�'A��1;K�R�&��t�8Rf�����4Q�d�}:f��;z݊^�"Q�~��)n�m<^�[e�A����Вu�B?Lș�`t��S�g�J[.��뱌��c�nQ����6���-f���OS��N�:�M�'v��On��|����JY�q�˕`3�$ډ�F�yJ��\�����
��_�b�^�m=�<u�zq��@X9R)���ϝ��v��&d1{W~��ĩɽ*Lu�y$�"{��Wis���y�|�(�(�Y�8Y��+�혯������n?aϳs!���)��_M�B�̺p]ZHڂ?,l��țn���@df�E�򥺕��0H�}N{α���/d&����*6�"/���6
�iK>bz�C�ʻ��[;IŅL�8cw��{�H\���HR�֭�cdƸ�ugg��ewWņ*E`��I�Nj�z� ��[��k�!m��1p�����Ԗ$��V)�
� ׍�(��%�������(�2}9�	I�
�.��Qp"�GH������.�����q:`�}{��ْ�l���$E�D�o��Fp��6K�]�6�m=Q2>X�P��?�Ű�3a-�5 1��(73r6J嘎��1V����ؼ)�c$K�\�D=���,�~�COr��[���hĝ@�B�$���,k^(�k@�|��7CRt��Ak㿫*,T��"������nQ��72uVw�wNR�����6]��Vb���X��m�6�g�V��Uku ��b6�����|�kj�o�a霩�Mˍ`��:�>�{.�L��+Fɝ�놸�Ҟu�L��e������c�z�ڛ8Fڪ�������>��Dh�lU�B^���0���m��{J�/�9qvx3���+Eb�qV�+�Q��
l��q_4�n60�d���K-�?1m�1����Q�ړٙ4-ښ��R[Z�ќQa��\I��5{I�9f5 ����~���5z�r���&����.8�O ��M:eTH废ž��*�����ڎ���*�V��)ꍌF,�������
�)8bx������8n��?�.��69�����5{}�O�K�,Ɍ��h���^�r��f��8|J8��r\�^��ri�u_�4q�>sw,��I�R�^��%<�W%�^��#%�7'-oޕ�i��Ji�gP�%(L����d�[�n�H��� _��iX�骪��9�b�`c�a���n7��t�%�q>q�p�/�-BTH������)3-�н7=������_��b���р0�(�4+����,n��|)�ۤƇ^^S'��*��qѶKإ���|~1Fsi��k�^�����T��Md�8rPO�[��n�n2O^ �d����R����x�u��bdʽ��|����fWg1܊���b]T�Gd�d�ƹb_~3��s@�X4#������*Z�>g������D�V�9��j����Y+�ѳ��!�p���7��ci���\w�~���[�]%��0e.H�hXРp�幹 ��/�B������.���j"qY�c@�lR/M��$.�����i�������y�#j�b$
>0�)K��aT��A��ǿ�r��b�� �)�͛p-���	�c��L����������iOM�n-M��� .jzv�H�Ż�O?>ɂ�槒�אe��$���l����c�G��6��np���KG����-f�,M8E���hW�V�zN9Xw$T���ѷX�b�&�5?���9�ˈ�\�qJ٤6�v|7����
�q��sܯ��	l��ZaRρ�w��������pvju�R%#���MQ
��r�ެ��'bۄ�IC�5VBɷԨ���s�� �lz��
뻡L��ؗ�������-5s��i`�"��޽z��5���
�r����T��y]�`.s�|�Q��
��&�M�3o�c]����o� 6����r�qW˝��=��*r�����O��2鋖��_�	Z�:b���W�_}�[g�~?xE�$��hWC',J:h9N�Uz��ݴ�ћ9y8��9��iB�\��`���o��$I��W�Fn��rp5�OT�-O�Г Ґ��=Lu>�C?E艀�g+�d�'��Nn�b&������#5
��NP�`?��A����^
$�*�Dc���'��B��%6p��jۗxӉ+�q��*�.E8�4���-^D�+�1���L0N�ʵ͐4�Tw`�_;���>y�t���$ ���#s�{�g����ӷ���Zw �N7eT�͞�
��U� ��]�X7��(��O���e�Eܞ<	qh� &<�߂�E���(�N�it:Gg�6��T
^C���+��������,x{k�hN��Z�����c����e�m�xc�;F���W�����Q�!��j1�Vc&�*W�>j�bB��	�I�E�c��=DnB�l��-�M���}U��s��s��S
�{�D����hW�"=Jo#� i&�r�0�V�u?���<R��"�t�p�9�#ů�o��7�:�����|y���<̓���9F�%�Ѧ+}X/��裯���o�Ȋ�6�]K'�/�����֮�I��HY�9�SD��He�j)oA�wXe�t�������:Y��,��������o;�î�aT��p�L=\V`��iUc��5I���
�M��Ĉ��w��=AL�n�E;*j�˵<�5G�jB�?~��PU|ϑG�[��"��wb�x�\�509&	=&q�m�qr}�u�L����qsk�4��Y�F�i�<�Κ���v�r��A�w)��≌�a�S��jJ���t|��j�i�P����Ye�k��Z�^~�=1��+?OrAm#��A;f:��Ic��7q��[����F&ںU�g�����W��~���v\xQG-��Z9e"0�W������x��
7|�Ʈ�n^fM��%���Q&�
4%&�@]L�v�-z֏��l(�_z��$�˴]h�A_���=.��7;{��^z�&e&����$�=��S��X��U���Л��ػ��,���c��e�'q��3P؄�7FO;������g\|`?��O;�JƠ�Ms���-�8p�``X�&�Д�p���v�^��׺ȱ�n�E�i-�u�(+�BԪ�(��֗:;c��O�}����-W�a�e�G�=��L&�����lc���_�Vx7E��+�&�>�
��ގ�����L��]��eZ�B	IZ�ۀ�&�Ծ�n]�ZY?�������{��w��D2ש��	@'�!ƧzI�5�=ay1�����o�x��6q�W*�'�>l�9y�(�3�P��5c���霨�k~]��'���R�
c:��6�e�ј��������ĐwiMAHX��]{_N�����|��!��&x�|���Z�{58O58�~1~�����)����68!�% -D�%N���E{p�J~��[�Ooڣ"C���p*�D�U���(�l:�/W�3>��փ�l��9��p�y`�G&�f�z��Q�(���-��*��Q�Tʺ�Zc�#��1g�I���"l0�k�C���,u�!Ƽ� ��g̝Z�r�J-�W���j�K����(A��u.�8#dud%�����bY�A}5e�C*l)�3��0������A�m����58�r�Em?����>I��	�9��<��g����J�gw�ꀭ�ńG�N5�FՔ1iDwsS4KQ�zc����21{�0�v��ş���B�^����k�,�b�´ҽ�7|��e(h�yU���Â}�����,Z��'�_��O^7�{(��=�$�y��0�^�N�͊M��}`�Î�~�TRv[&@�����6R������d���vf�E�hb$E����x�B�Z4���;�JTx捼mkhM;4��� �	�TN����:�{j��/�(j�gI�:�X	��7d�Y���L�~�_�*s/�v���rl*�g.���E�;n����]1�oT!�n�g�����
"�2vh�*�X�?���w<#�r�형�2����*����B��tp�F���~�����#����Әw7�)bn+�e�N�2��%���X{�D_׍#�!��i9�o�_k��.�/����L�U� ���%=�ĖU7� C~�M��VB�֦w	�/�<$*���a��2I��}�iV�����~ѥ%5+}�]��į_z<7�i�{00"K.c�ܬS�~��2і�p������#������"��6q�
�qH�>@�;P�V�HHh2�P�_ _�I�W6����XL����C�Y+C- ��uD���N�Ζ~y�h�2�`0��v[�p�,@��lG��5qr`�������QōY_)cb���������tQhE<��M	p�0���4Ê���sM�Y@��8�'2]&=,L?&ǣګ��\χ@w<JF�C46����!�{Z=��ϟ��%Q�C���W���s�e>�T�����8��â)�#�������L_p��M��Ct�_��=!1����\!��������h5���vVJ����#l:)�>�Q)���-w��8�("�]9��prK��W���h^J�so�s��d���k ���:=�� ���w���t��3m�gc}��h۩#&Y�O�����ŴSUj��Z����ja\ok�5sԶ��S��䷭�}i�-%5a�x_���\���T_5z�LTZU3����/�M%A	���Xѧ���^����Z"u�Zq`�T'[�hV^°m�x��>B%g;�؃T}:�2�K��_=#
@g���;���X�+Ӑ�4��j�!���7h�>ր��j�a�E�Df�R.�&�b���0�7��k���8�,�"�G^��چ��,���S���}f:L". T~��BI�����#�*ɣr�`�ؽˬ�qͨ�xxa��(�ݺ�n|�`�qϏ�x3�2Jv��2}&��
��f�:�_�j:#��N0���k����h�А-�d�����9{g��ک֎9ІP��
1�.ӽ�-�sH���m�G��OG��4
P��\�?�-d���H���5�]$
��Y�f�����M䵿(A�k����V��_Q+� Z��������X��a�����O=)ص����A\� /V�)vr(�&��̱'���o�dx��0~�G�y�6��
R��l٪�`����b�x+1�u�1���4_F�1TOm����a�c����ޑ�l �h.��(aF1|KO�L:�W�u<m��^�Aj�$��=�O�=D������L�U������T���P���3O�m� �ؤ�M��ޠ�]��������8����/�@Z.��a] [���rg��\
4��࿇F�����@��g�t�Ba(|ď����ϊerG�1�{������T��k��by��&
�*x\)4EdE���t:��h�J�Ǯ�8"��� �ױ@9� ����,Dd�.�'���з)�E������7�dV�n"��\L�<�8��p<.�u�@������CC��������4c>$kvx�b���4"D�Z���	#A�'Z��=�g��Z�+y��DJ����oƉ��~�1��"�Rg�P��*��ϒIA:��ETQ�}�	C�ێ�x0��������y��7ݜ�d��A`��jF]���\�f�j`"��4�=�����L�oLhDں̅���}`�	1���i��y���c��T�����FE9L2�1�)�P�7L��:�U�&�1!$[ �X�E���� �q~3ڿw�\�`�38'�	�P�m/�sx��gS�l�<������.�����WM4����:���u���:-Ȳߏ�?ܡ�^���Կ�q6��ޢ��ϩ_]IAh��=-5ϸcJav��X=h.ʬ�O0G]�<��u+��
Rɟ��"7y��FB̋��5����p��?��\o�3v��<+l.VL��wb���vo��lq��g��Ч�=�C��뵼@���d��8�XCD������%G�����3���?���u�QIc�[�WL�"1�	�jAa���e��a`��3KcM�����K� D�����,"�e��SD���� 5 � �0W��zfL�o{��F#X�2� �	�3gq���P�i���Z�\��kPsLA�+)N���섡�U3�M�*��^����us<z���҆N�@������P�#���	҈�T=9b��A�?R� nƁo���5=��*]��� ����f~�hRn�C	V(^t�ބKl����zK�^���v0�7�&���0}�mv��BFɮ�}Ӳ1�y����[�9f�.�=�)Azr(G<�f2�����(�`L�wwd�\���Jl�5�$���DVm)�,���	��D]�.�L�W����spkj�?в�jW���2�pD$�	�����M��3�`@,;C1��(3�H{94S�����ʹ����-r��b���3ݰl�u	@� ���
�� P���-�nT،j ���Zn�lrr"�z{7��RvofZ#�p�B�6�BT���b����o��,x���r��թe)`i���%�X5�Z:���i���n�C�NyZk�"X���Oh/<(�-��l��X3���u��<�:�޵��G�5Ĉ2D'0�Z� �=>X��j�A6��o6Y��:��r-�xI�'��{��R�=N�S`�F(�2�P�
Z-5�S��u�G�����������������"�z�)��U�4w]�ŀ�5�7�m����ߝ1!���(��͵6�x�P��y(��1�	U(&�J���ن(�f��0R�0��驤�}`V�Ή}W*�_�ܑ�}���jT�ۍU�?�ԥْ�����Vb3]���BÄ�Z���ݛԻ>���k;�ݤI�������t3�]r↖�[��������I�NE?��+�{��NY��,ի�APyP�N
98d��{�9ߖn��C�+�o�����D$p/azNQo�=�/
dȿ�h�fט�3�v��~2���q����1bi�~��u��ǿ����:��h�U@ɱ{V�-Ҟ��u��54sMénb܆�r�cZ��B�l �=�{��k���isE��8a}���U/�)H`�-��|S��W	���Mu�$���̟/����&g+�3<XV�6�P��+H�SMvbA���<�"v���)d���A��=~'Z1�h-5/+���F*����X��Ѓ�t�����<q��T!"�&q^��Û���[��1��^�;$��vH��d�_�'��n�8��s6�$=�{�H��Ǝ�EmP�I�肂@+h����- Mzl�^����imM�ۉ��y7��]��F�O���'�\�OV������[�V���j,6�]k���$�~�>�Qϸ*�{��L�j[ʜʿ�\~�*hڳ#�e��*�{|��#�+
9���� �h�X�v���/]��?�Y�i��A�j��O�>�W���^b+�e���8M��H�G ��]�0$<�Q-p��B,�E���؈�a�"�;�}�KgiMf��<���f�(�Q^CN�NGG�a����S���r҂�#G�i�(aUA-�za�X�f Y����j9,�c�j����W��u1+��G�)Z�g�y��k��A���)�.��ꑪm��GgZIV���_}�rB*��" �rB�S�`G����DV
�k2�<��1T�	���=�˷s����ID��98�Q`5�*����Dr�~r��iY|
?C~�/ݟ�&���H�6n���^��Zk\�O=@rx)�d�\q��Zl�F�`�!V��G�ڿ���ן�HO=<�`�Qui�r���'���=�����+�/�V��1F�v����+
�hOr��F�Q��~�x\ٰϗ��c���~q/()��^��r�[�lx�F��mG�gd0;	]"!�ܓw�]P��۬��^z�H��J����DEZ�����'�R���K��n��0)��6keJ���x70�A�_�6m@V�댬��h��!r�h�)��a48\g��/N 5�>/:3�6�~�"�GU�:�T)  �C�`rDd�/ߝ�<����+�us�*bn��ĵv`O<�ο*I}5�ֻ᫶��t�n�@�oj�T�rߣ��,;#ǽiE���Pq��a�����"y�/��8���e��!������7{uM�}� L9G!d*O��������wF��C������������M����({:����4N�0Jv�BV$���6O��󒪟n�<ێ���Z���q�nQ�����<ӏGǈlc��U8ɪ��*+���X���h�r��#���F��/�����$TF_�Pw�D���b��b�ZT@�q�'���i�?��c����Em<�@�K� ~$��뻸�����9��bdj=EUd�8Fr�<Z^D-���H��o�{e:�]��U%F˥mf��n-��,+g��v��®��p�U������V|iY �
�Ҥ����	 W0֤��n)F_6h�����C;��L+b�SC"��
+�/�T�/�~���*̢�
�IS]�!�C�U�t��7��J�l��A2�%oӿ?���P��֫�'T���+ORlbSI`��Q�ꌌZ�B[�F�����!�/�P�܂�&>��c����SU�.���;E]�~�
2EǺX�ؒ�l�!�.�ǯ��k*p�G�}�>�;�M����_��>�D���s{��K�">]\�A��������N��y<�.{�yLf
�|��l6;S�KH�7�� �^�A�XS>��(|����̚�;�_�ͨ��	n[@7�����B�'h.a�/��`�?�Ey,��B��յs���������ak�U�x%�3JRȽ�Ia��L������NmuY`)kȓb@>��S�є7嚖�[�B�$�����������n2�(�,ȫ��w�k��L��;��-�}ڒS�3ׁD.��ۀ`B	�;*'������$�Wjjo5d���	��2p��j��W��-8�Q!�[�v��c�p�
m��gz-��	�/tƘ盲�2�v�V�� �<�8�nt� �J;��s:��ۿk/c�~���n�O�o�ͳ���d�Ǣ�m�^Zs%�/(g�Ơ�sY�/iZ*o�IuG0JE���������CݴYS/�|ߒ����\8��кS�NX=�>g�[zOfC�	��D1z�����` ~���|ĹB�Xb%�V�j:��nI�h��|�!5��
�����o�$�h����ox_�/� �L܇b|��ݿ��bbM!6��Vc-7���Ŋ���h����;v�#���g�mǚ�E��!OŐ����j;������;�^�-⇮}@�C"t5����/I�������;�}��*L��_p�6�쪫d��mć���]ƾ� �[ed[�������ة�6X�#��Pn.@�Y���ć��ŵ��E@��*��.�	�NM��]cv"�F0�G��]h��0��?�U
�.X_���X����W�>��)��h�,��ݚK� �;3�<2�Y��[��l����Y��e�Ă\�¤3�j�SM�}�^��P����r�!�MM�.���F��G�{Dh^�\E�	��4�Y�&n�����)�gT0dj����d2>D���������]o��]��z�)'#L���(��+T=�wF�)�rX�5s�[��y^�=��˷ckIz���JU�d_ �~@�Jybd��H�Ө6��x��Z�x���yW1�\*ኽ�T��v�@���ES�)2��(���W��KY�9�:d/#�0�` �a~b�+�YG;f��k'j�>ܧ*	0��v��|<��q[���I��0)a)�ʳ<�(�A���O�nQWp?�L�EۣDWdd 
:�׼��璞�3�R���S*eK�v��T�1o�>�I��ɂ�ɯ�"�����֣���'Ҷ�5c�R��o(�w�8�K����RƎ��9��Ԑ9��8C��1
���B��J��o�21
�9�v�X�#�lA�XS����H�(;?��3n%���Ly�#&kf.�^z�j~���.g�	����~��4N'��E�lo����(<��`5��&yɪtq#��D���iy�1&w�}�2�ze5Έ!V�6��	��Z���E���E�9��А�%���5�D�Y3e�W
�7�%Jq�M�m�@��82`�c�Y�Kw��P���3u[1Z�a�;�*a��ܵ�9���=��dD;��11��)5�*J¢��k���S���d�<h�cEA��6�j�-����$�{.C�.P=rE��������REn��2�)�[�����"�o� ��8p21�؟\�������"+��fG�vQ�2�$ņ����Ҕ��6���Y���r��6wV���􅕆�7t���C�8h���=$y��/�,,��)nW�T��W�cs�zO��΢�V�f��<�T�B�7EgJcB��~���F5�g��vة�v�+�zb��s�Y�6��O[������FqwN�o���=*��G������Q{�O���T�����<P��Uiw71���l�|��-���E�����Vq��V�����`�e��R��TUp�x�ۊ��z~�P�8cu=q�U�w%J��]��D�Ȩ�9�,$m�1����e�(Wg�ԧ�`n&IfϠ�w��p��0D���T�<\Zr=�P��X6��I�M�_:u1�@��&���8��v�D�M%�Č��N6�:���%��6L�<��):��S@�Y`ό���!4,�؇A�� W)Nn�N�O�j?��|d#A��eSș`��ug ����i�%�0O
:��i�����V����M���//Iq��D�Z����}�K�	�̸c��+*�t>��t\cb�NΜ�Lf�k�|��<V�? �8���|213&���
U��`p�� ��)^ݜ���]"wб��^EH�h<hv��u�}��7N�c�_�D��&y�Q�}�""B��!��F�vHv@�e�?`����y��b��y'���F�C�t��a�cu"�8�!�R)�B���e��W��?�	�⏱Ɠ�S���jv���>{(��ey���ה�k�8D�.d.q�-U�~���7;`��*�Kf]{����.�9Ư�K�`m0��r�v4�E@(b�s:��[�@��gg�J�G1K���<7v]X���u�����%�Λ��������]`�W`_��F1T����@�S�=�ߕA�L81nvg�_'$��e|�5��-q���1"Sj�3�!#�����uдj��Ǿ�w?�0%�Io����=ĭh��_�c�;�U�C�babt�o90V!�q��Y���:��c�\ �A���Q��x����e��~�`7.�<s߅*r'O9[�E�.�Kӷ�:n8坢
�?��0d8o���L�P��xe(�X�P�`2˲�`���9m�s�(^ߔr��=��MC���)$!�pv�D��x��� ��;��h萐��sګ6�f6�y�;~�I"��%��[������^DW,CI:��^�=�J��������@L���+�x����o�a7ϥ�F��x�,�a����<��Gǥ�;��ِ��T���>���!1���C�}J���T^.� Y���!��+}�#�jQx�JD<� ����5��=�Im�F�~�� ͘��Ո[�_��e�+Y,��R,���wZ��tH�}�ճ��/ﵲ�c���.óm�%�`}�9�7��!�_���g`�����ݖ%}kb �(�<v�j�Zg��9�.�ǧ!�QS�b:�/���zl���$�2%�m����8H�A.Yx��k.23�`�*������rb���W;@�}'�����\�(p��@�H���x�+�_�|�ce�QT_��S�E�h���\����1L2�T���N��^�.�O�t��f�p�4�輠�W�����h"Q�|R73��t[}�"ϔ�ȠԋG�t�]89��<���P@�N�(��&O�����?�j���! Q�̡����=�U��F�-%�0��� ���w.a_�.�1MO������N�X�zq-��n�2�� }=��>� ���h�z�l���*c�
��!�&���8�J��1�33=Y!���O��C�v1���f�Q��.	&�|���̽X<���ƣ�s�}���x�_�r�	�wR��E\��Q9�]��}�P�DC�	zwL+"�s.�,i��WB?x:�P�+G�"�K�ǩ�=G���6��w� .#��T�^�b��+�P{f�$)����������!���o>Kq����K\��z7�;��-���=#�?^���6`b����`��ܲ�p-$��4���F���;����t�,M�4�}�����fe�hSu�`P�5�?��@��$=媊9�#�^�Ǆ�tc82x,�=U���%Iqo�y �SM��Hp,D��d�w7������S9�~,� T�9�Ed)���Np�I/���%�[�C`A�1[UI�m��)S��i��z���� �s�8j��}���$1�7���u�GTIE��O�u�ކz����ڛ���I��m���k(�QH��x����v�O�x�5
�f�[Y�|	�J6�!�tv���3��E	ʂB��O"I
�&9'>�S�C���E� ���T���]�}X�Ӌ�a�g�6�q`�������רn)��έP��l��F�_
.J|�S�S3Boȫ�<Ŭ�Q�w��B���c�Q,����P�@�A�����Zef[qsJQ��u&��B���/�aPF~h<	���iD�`��Ac���f'^��ɐ��挊�.����N�V��˦*<�7�ŭu'1 ���~�^���NA����Hpc��tտ�0���e�E=Ð=
�{_4	KPrsޯm���g����,G2�W��)�b�9c���ݵ��Hg�?�<�nV]ztl�	+IWx*o���l�8�w
�.v(z��n��� ����\�0éP�U��6,����������_ߩ�AZ�����0��bYEL���c@j���>��C��ȼ��tܛ��b&�5�Zt���ԥt����b��-��8��qɸ|�*��A���ޝ�ۺ���^%c�rbN�4��AP"_T�� �E$�u��G��0��Ȃ)���X�}�6� ��L�� w��i��3��"ڀ�/re�������x��c���J`藧�'�]��1��~rN��a:�8��#�X�pl�����ĺ	�����}�=5ra�C�qn�@'�����-Q�Zh[�,�_���!��4Ud�^�`/�N||Vo-���qȥ�� �p��!���ڻ�1r��q2������H�@��P���"FAǮ&��*C3�J��jh�o��BUU��b�G �����2,wB�oh����@��:2�2�ߓ��V� ;C;~!�bъ�s~�K/�w�� g��!d�Vpc�j��S�T"϶�����sů��i4>�dҊ$=������_�]��(�м�7���|F��u��b�9������-jizow��-Ɖ���w����q��,�Є�$�؀ٳ%m�n��~דGQ�r�4z�����2��&�+�"{��3����]V&m�f��X���$�n�u�;.���ϼ�Ȥ�&��8�7;�i�D*��~á�t�Z��z��K��-�듾���|yu@]p�k2E|8�uO����5`��Xo _FNw�I�'��-�'�-����6^��
���~�G쳾�G���k� r�ݒ 5��#�Bf�\����j�#�Ϫ�5��K�v���OGK)�$���O���\.�uP#A�3���Wǯ�_-�_�ݥ����2�Ӏ���X���w>�/��a�_Y��q�IE�!���\F��ֆEKCA�%��E8)����y�|iT�v�,�E�j�u΁�4������R��tUj���\���V����O��,2(����G����t�3l�����H�!���ɫݴjn��X�hy@�d5C�F�Nv�PfQ�SQ-�t!/ �d8�vf~$	�&��	��f�~��0�r^�ረĹ�&��/be�6R�1���r��g��J[��d�R���?��b��ʝ�U*�_����6�@�H`��x�7桘�GA���O�у�̨�i�)h☋�Zn[!�� !sIo!YvtBeb�#�8;�],�f�~h��k�4^P͒�.����>+�֣�6��^���cUHU:��1�ރS� g�Q��hȊ�����Q)��w��i�*��{�[k1>7�+�C���f
��V
�Ğ21�
$
j0�2'T*�v��%�ʖ�6G4�?7��e�	��~�I��"����e�5�X�Ll��x:m�u>�����n�Sǰ%z#���x�����n����c	j} 
�Zo<`�)N<]�_A]�<A�5U��Epy��r��4��p.���ؘ	���_L1��3�� �ѫ�e�������s�� ��K��؊�!���B�s)��ả� ��9��!oM����6B>bӵ�%:u�<���y�������+i�{��S��1����O�V��U�����Ϛ	�`�D���X�a�J�8��2(k���2̒&%.�<��FEM��6v���Y:(G�.� 	��G�1c��Lv�T)>,F�|��T�;ocm���}�Л+ʭq�aN/b���H�d�3���v��K�nzE�+^�mS�҉+�S�@s	�d��f�8��8LZ��⨜r��s���E���-��>��(c��ȉ(����̡���-=�#���n}@�F<���v�C�F&��*�6���V�ޢ��Ώ�酸C����Y���Ԡ��:Gs��jPm���XTH�`ۯ���B�ThX'"�RI���p���W���(a�򚝫��RI`���b��� 3�nP�o)�ƻ���SJQ�kb9C���| ac��(��1fWl<mv1�I +���y \��,�g�欯��;��.�YƜ HB��^W.�2�;#?�}O�R
a��(+X�J�w��<l�W�Z�v��j�:ޤ0 %Ǆ}I!��V��?z+�D�1��a��V�1ĕ�B��B�x~�lk.EH[�ǜ^����O=�2G�K7GlV�����Z����z�6�/.mB��.�����K���� �ܘSe�F�%<��h��,UQ^c�Ax��_f���wD`C�����=*�u��z+����/��Ĳ�\�O9�p����~�� �ywE�Ӽp&�O��B%#N_}Z�XK���q(��U�Q/A��W�+7 #�d������`��S� Bߕ��ڋrY�]�����.�6��tC����wt�&f�޽/��'���RӞD��G}s%�)P1;E�������F�qB���"\�����7���
���zorb��A[r�,W��������~�4q��+$D�ں�{��q���J�������g=�S��-1���-#�$�6�H��$�j.��ڙ{��%׾��ܵx�^���&�nX�w�ݨĞ�[&+,����g����t�4�#�������6�rq��IX�0	ʹH.�Y�V�c`H�#�<;���x�n�mP/�^B�1��K�;�K�����'8/�k��ZL�����D#�S
��E$d�T��h���Y��U�ܱ�ұOT�^��?*��EF�= ��a��@s�M�숧P�Կ�Ԑ��W���� �^�J��:��
�G0Kz�P�B�c�E�H����?���[՗W�5�1a��]��Mc���\����"Ҡ(I�q|�����vQR��rʯ }޷�j<>=�^1Yiʚ����|��ю�\6���z����,��!u(�w�)ﲹ�v�Hve�)����✷��g2o��g���'B�U*�p�%�����-;�ձE��V��8GV=*��>V��@�
�C�����I�Q6L꯯�Ǡ`;����|C���5��i4�����r�����e�Z���O�
eh�/������0;�e��݈�K��sL����rv�'�����o��a�z�A���Tp�G@�P�[�%���4�FV��zY#�Ƽ�G7*6��DO�1r��N%5܈z�8���'F��7�\��aն4l��'Lt}�&{}=�9�����˚߶�b��Ċ@H'SN,�������$��sP8��E�?!�ޝ#G�l��΅�(;i�/]�k�rq��~��؂Y*F�WJ�~e��I�>��2[�s7[�梇0v��	E_	��z�m�T��Zq�1��H��+�ݠl�7kD��>j.W9�ѯ���SG�3��F�\%�\]�ȓ0-'qԃ7�4�@%dI9TӃ��'Ȣ�fw�mڒW�&_m������~r�ze���t-	�!��1^��񭂶8G6̼��{��[?�o�%�g:ʬ���Q����d�F�ay�G���>��D�\N,yƴɒJ��xL�
�7|��M߻�"}ڡ�O�J��y����v�s�x�hx���S*6�$N6N������hy�X���g�l��YG�����wӏ����2��aC����P"m���"�2l��0t����L	�4�E�>�� %ķG*�d��2 ȧ���(�3��$��=���#�M�1y�B�E��.}���a�-���k�EF&7�Bj}"`�R�s�b��-ԁyh���C�ku��zZY��mx ����l�Fٵ��C����J�����S%�'еi��ў�h[>;����FY��4����KwlTÈ)��&�Gű��v+Ar��N�c���'RB�<,x�w�\[���qDK��˞�k����v�n��Y�My�͇��<KT+�Q���B�,Vwp�e�<nz֛�Y�y����m, G�6�;���%��pp���X]��rB�L��d��n�����C��?��$�z�|y7ƙjl=��H�'�W4��u�v<Jz��H'e�w"��io�pr���1��viy"�=�����	�1��5SRVM*��g�����Y���n����U=�mz,�W��3�CBM���uv���聗.�7�LL�3MY��gH�V�x�@�*�b V���&���	eލ�!�8�sG�N��V�2��Ik�������H
�B����	;�7 ��&P?�_��U�.���jw��8�Uu3��P�jd�`O�3�ڛ�!#�eҌZֻ:����� ���S�h�x%��ދe�~�n�ڡ~��:��T�/`m�fe!z��O�3�bZZ�1]7��$.#/b��㍩[�Z%c/U�.�Q9*�	���8��",Tn&�=�7��]��q���)�U�B&d!+fԌ+�iP=����+T،��G#���6�&�߭��Qտ�e��pz9��-�R����~�M}�,AĈ�W��$h�/*g3�:����19x(`4���2�� � ן��x;8�(��gٲ�\[V��ڙ T%��*�4�����(E�h^H+ќa���
vQ~8W�X�5�(��SW�x�B��z��
*Vg!U�db�^D��u� ����E���ft��i��wۜ`�d����2� �wOr�%�_�����z��x�#��G�ʁ�kKR�S��š�y�O�����>�����:��U;���ҳ��|� ;��
�'���1�J+��2�2f'qV�L������x��?�qLQbd���η�C���f$W��ڏ$������~
C�`'3YJȉa��-i0�v9j��Id:P��S�J��$^�/U�e�rI� ������ :K�x�P������e��}	�:}�b�k�qw�R�x�j�v�A>/����A�[rJ���������ĶQ��
F˔Ċ>���'>�ֲ�;y�k��˙5��{d����{|�
��a4���ы�Cm�J��`���w><�b�Q��kK�w�r����?��zz�d!�@�|�r3oӼ�*��֨�Es�����������S�T�F}�kgР���9q����M�V㲝}�h��ķ�G��ى��mU�|����i��i����<�)��S\ٕ��rZ��޻��M����-��bK&��Y�B�*�.�\�i/˦GV�1U�,̎Z�H�ξ�����S�sƚ��;���k�]���c[(�OI<��_�dO `+�,�*��h!��*e^��Cj��{f��@wc���gn�����饮OA��!��� ��wa���jv��"�h铍t3S[�UZ��Zb���Kp)eoь�Y!���hL�g�L1��@����a-�V��`���'���M�q����A�=L�"�;�y{���P�ud�sL1z
(��2a�c�d��lp������3�L1����H�l������d��%���6�ە�zvj"�"PlPʖ?�*�I����{9�{x���K��� nv��uQs�*���b�qiJ\֘P�T|���Bo�~};d��i6�FL<���H�)s����G����Y}���������<��G��})&./n$��yO��ol��5�a�#���y��j⢮�wM��@��7N"
��G�[C����U�>��D��>�{
����d@�-��&]ҧ+�n�����W������4$�?u��IE~�/|��#H؂�z�v.�:��MOǉwz��,=	�x��|���P�J��x����)��_�kյ%T�;����5%�M���(�8��)���[��US��A�+�^%w:|��_�A�딸~�^�-�¥�� �
4� �FzI4�{ ���=j n�C��cs����{�o��&;E�����8����.�}XH;ЊO�goB���>^q��ԭ'ǁ��Q)@\ܖ�k���*��p^d���*(���Նgjo��1u�\�ڻ��[������~��{"�G_-�/[y���'۽P"h'u6ȣ��W���t�9�����@�.U�P������d�9�rk��&]_*���'�exRہa�gn�4���C(+�e�s������bJ�B���]��1)l#`h�궞h�)$��zhxR�.P�wIhU����Q�uI��Z� ���#�D��-z�X���#�C:�H���=r ��b߈V��8��';Su�Y��0�}uI�"$�}��s5<�����
���
�Ņ�Z�Af$'�I��G�|d �N#�Q��	�^���=�mf��ˑVŇۄ�7�_L>�ٓJ80��'�7	%R�9��(E��`l���� �'�8�M׭�ƭ�B5-���.B���sx�*�M�p���0sI����G$�#�1�$�F6H�B"�ܟ�$�ܼ�'�UA��F��g	{ة{��6���S���5�w�E��(<7�'��� k�	�\j\��������Q�����a�?��?O�P�~#����<҅�����ɮ�Y�
 �6z����b�:���e��yE_��9��L-�M)�ַ��:��,�Ǧ��¼��V���cA�ڢ��፬Rm��jm���aK,�LL����x�2�V�fF�RÊo�M�p�!�GF�Qy����_Gh�v�N�3���_�O�g3�9��7%�k��+�։I��c�>�&�7:�[����iz��7�&u���z@ԟ��ev�]F�>�(і"g��8蔶` O_�m�9Ua�����$
�OU���mK�)K&�,�@�`s��6���Y���9����j2ZNB�
<�����M@x�w�� �(��* ���%�y�KTXd0��?\�\^)�۝����6N��^!����%����>�8�}���\����u�ߴn�{4(?��.��̠���E�6Ϊ�L�\��[�����DSt#Ю���v��}��O|��o#C��x��/J��3S�˙@�*�VUP�=־aK�#KT�%����ָ٢��g��䂸·����i!�n
=�z��ק�em>C#����t���upbt�Ҹ�Z���]Ĵ�j;��1H3ؼ�|d{D%�A� ��3�aU�;~��(�V�E̎�M�ޭ�N�^�hyS'��-%#
x��ʢ�^[�v)�Í|��gFr�r1��ﰁ�5LO��?��/T��A�&��t�2�n�;W����	�@�ϫ�Su|�lb�=#���?��>�"�D��"��a�>-�Ė��Z����	�T��d�h���s"��_��enq��ce��45K��uS0+�QFf&R�SS����m[�+��_*4�ge٤J_
Q�O!�`��47�)�F'2��8LŨ��A�[�C!f�~:n�i��0��������_��MQ��#�2����vkS)	,DMS.e�Y����Ϣ�����$����鈓�[�����t���X`��������Tt��v��t?�R�{]��n*>۳����Ⱥ���?M擣4>�7�@f�bL�ݬl�����Q��!���=|��`7�>x*�G��WJ� �8��jRr�,��N��s���C9�t?��<钴2���;�[����s����k?��3}<A�_�\��K�	��Q����.����d'ڮL��k%o��������`����2T�>�bf?�?��ρ��xX�ߣ���?)�[�X.16M��W�JI��Ⱞ9g�rM��/�N{VQ���\�'�zĺ�g�Ϊ��dǲ���� 9㹢?@/n�����C�&�[�?_�r𵧫Ț΢��L2��4MT���n���H
�?0�}��Ϋ�D):[�v�-��S!ArϿ�9�rTg�LR܏wLb<�ϗ��&�6^ŗ���,OnF�q\i�1�r��'Nj��