-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ur1gYNPexbqkEIJEYS/DrJmB+YFOD4S3dzhObPRn2nRgbRmTlMG1IRM6k7k+5mlS/2iixdBEk9Ib
7yS0vvWCJD5vHEaijbD7KOrCh0rSESmZZlEVbF9+4z+lrQESPeRRtWJSmlOEmVP9J1FWJPwevbFG
xEdFU+tCcOYyYDBlJkgN7hNhVnGuY2+XcMtjNS2YUhfr3Cyqoq775qCM2deb/AFiCy7nFeyx4PBJ
usFSRhXb9uJA0P+IsgtXGU0/xntfX+bFfTVYXl0i5rrVjqqcLKCj3D7mJFKkJX9rUhL4Ib82+aeI
ToDNOZLOZ+9Cn9wCHZIxAUWc9xng9jUpN1hQUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13936)
`protect data_block
ndfOXN3W9yrpswgIpM+wOd/oi3uDVtSxbLORoMcXSL2Aa6pJIZDk1uvFsSN8ro7sIUyUimWUeAms
EfaMOxY1qS8AF8IBW3QxOd4Lwqzh2in311n6O5pxgHKHtZ35Apuw+9j5Kbtgvk5seYd0shmEBgwi
wfGGLCj+e4LkfpOxKI97u+JdcYpu3iLMG9eajSVUuKL3ykPGcZ0UGJIf++mj0u4r7G4hBrF2jzbm
+qOyVn6/bAP/7LFCp9VDXJNNqijE2N2Ckq5eTD4er6+35NObE+SdpwryExzn9dyDkApmDO6s/wC9
mU1V7Y9Pv76ggh65JFq06uTfZ9P3gh3FXEPON05kmVNcT4IsB1V2dZF/wAyPrarXyTlkQDHOhrjs
ZCWMIc2Ka5fC0pZ8Ly3Vc9C+93fW0C44DxE1SbRD5lCjGR2UxRUeMMNCBMEVU0maAkTV1dlVayiL
xJdQtyUhTSh5pzh5Z0QFyzT3QVwxkbJ4MFbbJbcTfBuD2Dpr6rhNoKztZ/wUTBFrs0iV9g/69R97
NuWjq1TMYvqPJAlF93Mu5UQbhedf938L2pV3LAfb3vK3wgqg3OE/FNfBgpT61kVNudqu3L6aIrDH
AlyiHmQE1yhvLbQtk1Hqi0hqYiEC0RDF/8vfNvZ00cPkE7Mz2lg+Rxz4/yrQZBRxNKNPF+SGHoE/
Sdpc82XiqRyFxNxYMDupTYAdOaLjAirfawD5BKbrRs1dAYf21iK6fDPs+tU32SPMUyo3qmkp3Zv2
azsdKizOkSgtMXoUyxx8UkF8ggKJ50/qJGGJipmTfpXlXXbEwK27sB057I32wE9I7CCqXFfKm+N9
IGdIJgbHklO4dBY2vBJHRg2Aau3hb6Hq0wL+3QAnMVBlsW6C9YPD8Xor5798mnJiXDuUE6XVbXP2
kCHgNLvqktVo3GiDOwY29bTqJdocpvOtIlzcANls6Scq1aHLCsxsvIWqW1IbexkL4roZI26l39qT
F1lCnbjMRSDtgmXR4DHrKAZ62JPP4cFHmNkaqnlj0Z7gHoOufDFLm3hnfYiP2NG6U1C8OR+yul5P
kiMg9YBAYMD+uvbFWzk9EH4xrw2DFukOyf5YecRKNbM0AHSclX/F1toOYgqHoL2nwbUjJPsroKgD
opv7dsfBEGcez+/KdGPJAnaV1hdEvUJUmOPnJbtFGu8maF6oP7gz9q487V3BtJr191jW41wCikRe
HVR/sYrYdZlpz93UqdfsLXNzT0GM6SrxQhtqtIKHOTgQii/oKFhZw6KP4hX4/ShYqLWKKX62UiQD
F1+akfF6DUUTiX1xV7KvqDIIJXw3N3E1DuiYM+4eYBpdRv51J5KRAyZQl6p2f3NI3m23U0mKgs3G
DAb6okFhlTFEa8J2pcCm3u4BmiXiwaTjD0K9nEcgI12JrjFvicz1NIP6Bfy6JljOt1STyroFetrE
by7QCqddoEIzBOiK+hyX6LB/qC9TvMfzAwFarnImr52YQtR9eAMR5rPpzKPCFTgKj/wduUH3dZqZ
NDwxk0wUiwOxNtTdbs+I+v3fwS8HOHlbQMxVWl+NemB8BNUTGcyLCDUnnTLsWQHtu4fVSDbCI6l0
XEnsJmEhweAUlgklBRGgi+jBB1Ev8hif/xe7blj2Rafvy3MZWwINUSk5tsWBg99vP0K7ScAZuhxY
qPllUYxsecwCUlehKF72kdTcYcRYyhCs2nRaYdyu+Rn5ci5HeiVDgeCmq8yY2GhlC++WqWnLAzIB
C6C4RFl4Vts8/qP8TpFAsspCvmKCYSl0Ks3nApMxikwb9SwlGi20bzPp15O+fGZRB5+wlywA2hIb
kF3eKbPdNmAUyV+niaCXv20e+i5gH9s4VbUUlT02eeEGXnvlsJGLM6Az7QcX0kVLMfZglGYo2kg9
rBBOXFxSNSiQAeqhgpxoTN4dtxShViT5iaoH1T4Cic8oP8iNON8lKsX1QKJopW4FnZDe5bjdj7/W
MgA0yHQhVWG8LGcvVTBwTUhl5jrWQawLzwelOVGBea6MWFhCFj4fRccGIwzFPzb/hmHUilz0i1j+
IS+p0gGMXQy/Olk8xX6c7wiKgdCRO5WnXF170eacuFhFFrZyTi0HTpT67HcFlDGDXUHhFVqSCBHj
qwmen3R6RrWeQMobdq17veUiMJAKwpBlJqLpfDpYYCQ2eFuzWiWi/hbSGD5obOCVt4QrPh12FzgR
/yq+YNGkkArvZcyH3uOWAwAQlUQpJ7Tdn0Czbp6FVBfvYxFqcPUKBK8sZMO9xd3JfECiSp8r5sQ6
OWgknxpSYd6ncTkPA+F//9ehFFHYOnkZ8gQSx3M8jsI93zR1jc5CdpX6I1IjN3d5x+NUQwwkjea9
TLX8Kq3Vs+M+6UJrdbFaqDykFjswQMFd8KcFDbCzYSdDJwupXTULYIf7lGhs0dDBlWOQbEQkek9e
zA0DkoO81EMLdOWXiLE6dDqOKBZngyr9Nx63JZffyX4ycOIemqlLxvPtyx0RqN3ZMXb2lPQL1OHB
GRXkJbgLf19IY3BcvwgwWx+T4YcTFOMXOqXP8XW+0qIkIjfQs0qwYutFLW5V0UnFwHujmqFkI8cV
h3VvCl8O8nsmjeLVMaGzBC7EJKtFxkf6sOj6u1Fk+zrqU94bwGgWlNN6nKnC5BO2AfOIWUNlmOO3
84JwXgCcsF0tL0ixurd/23rh3TqfE7TqJv3GoXXSNmT1E1T+q7SJaLv7rJi1/4plHdh+N3XVghwb
2SGaHTZTuH89vo1HU39aC+MdeFMg+KdLVNeDyDN4DapG9lJKkUvuuL904dk8ae3cg/9VEp1RSEs6
Gne+GC4yokhpYVBSozk+pdLVuXQY/9GuGA2nF1atlAiI3RcfvnvRlYEDvY9CFeMLPZg6MF4Pl0TH
wdPuBOhsgxxtwBbua7DXz+LryDmVP1NuInHAdXbobtVvwT5dPiQR/fWdbr4y1MhM3otkNgwYzp59
L8zfLyJ/Nev2lzsr/i+uZYz0lXKiyUPU0BfeuOXCaJ9ujYeWZUlmUDdqfMpcjQZZrbrKTYB53+YP
95cOiOxcdbimup5IMBOGbX/B50VDoAWAy1mFXymIWfNFBAZwmQe9OL/vHSWJFmfwyyJw2qDSqjEn
rkbDxAY6izstISKbZWxtGpXaWJOsF49Sj1oGBV1YvYbugFFYhdmy7XVSvI3O6T9GwXHn9imCxzGG
ao925/Wr228vD0i1xRI3kK0UblKkKvMNg/EI7cmJ4RaIQlPLf/jTWyIl1WBhxplHKQoR8vq+sEqh
hzHTRfj/u4MlzuDLGoVIZzYDTv2PnAB6Xv8NAEUMUvN5vM3iTqZfAzhIQf+tHR3xySCia8OyhMhg
Qatj6qhkLIOlyJPr5kfdQJPdJlCLdjs6ZVqm75wpBKh2/5nDcuT34SNxpa4Jawj7QKzP5spaoRfC
PHbWG86LPsK0I4mVGNhDtDCqvsh+IMKk3p++D6BpecsHUIXvRhIdYkWP3ufl03SzLWSb/jy6KFT6
hR9Qiht3hKb50NcqbCqtkBSSMiF8UhI6vnABhaX2liWeFamYSpVC+7PQo4EoG4XZ7P0n2Rd3e6ar
2JQ1dfXIz3CbPZJla0fJfLq2ukyJ+fqLv7cpDMV00y9huN+GfEYdgz6c59vKvLM5gbgVVHTqkv9A
hTz3Ex9H+fxMHDUkgSxxXPXpTekcTeE5lTUofHfB9W+uqQdSrolYlzJVN7zQFCrec9aukPhkPLQJ
k2ArHw41kiCzHegQFVE81Hlox8DF1tKlbp/Gq5ipWCWhLtkvnuxAOHFrcmyEV0NFTqNWw4VUQB3b
c/jWg3HU/r3vSal+fb4ZsRUG+LWYaPM03xusotuhJHfYOG66UgxpFrIWXQ/yV70WaCIwZJGu/LkV
UmRm2zh905EzYQSVSlu6xLPpTQKY13t/m45f0/5tSLctb2yQ13xWj2sJ3zfi4tusIX4Npr6lzBN4
5+NgcGVRyDYzcx7PsIfuTTq5m/5VK1hqPnfdrbOJ3DPdRiQYjhZbn2Siftfp7JSBeGd9oJAIHCeB
bCz6CJvcySpaWeP/k9mPMbRx4KGuzX5sG0AYwdZqouIUV5yj5auoONNJhy18na58WdzwD8cAb0Nf
ZaGZymgqplTfEW350+f71XM60t+9e5iMtTWyQQ7HJE6Ia6kI8pTR+QDFSd6oHmz+JmExK0DeHeUv
VF3hsWMzw2jrN6H4lA83C4zezd9Ybphv/x06whSr7r/8KwQGfDbeGDPLkvBAlbsJXGTO121VaTdx
gqQXJIiouOYOLVkVXqV6YJoZ+rqqGbUd03dMHvP8QlPo6RPZrgpHt35T1AHymL83oac7l9T1Qpt/
yVTWQnCBbL0uB6wlXUh5V6aRqZgYLYVJkkBf9toIKjzaGoTZtUI5T6qRcfYztF7Zv5UQE6dQYLdj
IA8y2ptqyzg5Q0++BFh3GzM+f8UIR6k5UnIFEzEierWrGpfGMGgEAfcw/7r8hJE4VKWxtJNxzNBP
AMTmCT+ww21xMxkbZgS+xVXzIpWy7PYKOgRGay+OKuops7g15cz7vLZ+UlmWlCOO45/qsrMYAiB0
id74ti/1IeZxyPDu6RjXNVXcYV7yWWHr4p8Wxp9lid/2Dqb3OmOA9VarohMEQiLWF7dQpSBtwlb+
XvouK+AAbVhgopC76JI7DM6s7K/OAL3Gx4grpPMSgsRqnh+spqW7mm/2fO3mJaSNJ39O2cNmme1J
lmoacILHHYrOlK162CGc56wosb762sO2C4MXSYhTRE+Mq7WKXy94J5iZ/3+hKYFcq8vguD6TU6ul
91yo/L4sk3ypucoIqLd3etBMCrSeZwByebCX6PFyCx4exjMYx65uFtc2nhqZrcSEYUVNOiCCmWk/
yoffH2ItI4t/kgl2+ZBCAxJCKKsCAOxzMSkFDx8j2B9lTuAem3Y0Q77+e95y2rOECIjU6ejUQZBm
35JgWfDibHg7EU/OnczH7pc0lCSvEuwWTTCAssuMvH44msH1oAEG8uoQMIH5+DqCCTHDJu+uh/CY
c0P9fR3k8yDKnfdjVBph2k+ztFAZ6HDsAoaYUpdhUjwKBbpgzU6UPBwN8Idoof/7wJ7O/ZqlNPHZ
PtmmHrcME3w+QgNM66FUZagfs/s9Ap9a7jD6EJ5ZkrllPjgVa8wlb7QaVB29fS39kIzCspUMZOlC
kDJGIzsACdNGyaKmpVnwi2acWgLX0d2cG1elrbHmDCoXAbN5X6U3x0INh0SIsvNPlBAPX0bn9m0c
gz+i5cxVPLNJhk9Wga7fujwWJAxSZi5kUTI1+1RdD7jOVqG5DSasmQIhCeOSTXyqvrzK1nYAwcwB
DTCiKFW69hTqlAN85kHvDutxjpxiE1ZX/Rv2tYrX9WlvagfvLV4MbIsGe+Edj3XjGUD3H7pzFCMG
Cb8Sqoe26am/z3Mg1MkNrK0KEpB0BN3Aq0N2U2MT4ZVxV/BiMUPuhOXKdbwe1JlTJgEUGNoxBvAe
lAm0kxiXt+OcwTxLnd66TdKTmpeapuDOJ696emYpbhIRRhiERBhOr5AvKuTMUdcKFvBIlsfR3oEq
GI1HHwDPNZNMNl5aI3ajcekKMHwhiBINgKLIsN3e5Py+W+N1uk8F3k8vxQ0rQ5w+u8ZV65xLLZts
u/Ts77e+SzYOawBtZDe4yKjS04I3/ignAfcBdLaQAFOBcRWGvG1yNmr6QPbXx2jQWC1wALaWkkIV
z7pTsbfIZ0ywyHi50kAIR3dnvpdHR2cEuz8cRxysKZ2admJn7qofXRFrgdwReZD8cvUzqiGHa459
qv4Ox9ujfkuc/DrdDrrN7bucdFtFLq3F8uyZWIOeR728PRXiRLu2ZpUsJ5VTNBAUqxhyJxidRvY0
HVBmkwIBvEn/W15tB2GNMVfXPSMG6wUMZvnMvcTxCL6KQNE7xx2PQoX1u3NU0HT4xIKcS16YJZiJ
EfZpnILwnu2tlreDzeta4NUiGLzgoDdSCoI+Rnmdaun7f7FH+1XjgIPSxVRWJgeFF+ZbO5BJMw2U
ql5RQJt8NYl4NN7d1ShfJue5XvtVV+6/5M4cOhgzGWYIjeBlAIsT3nHLqBR4EQaC7zps2O/E60Sr
dT/NuBfUHo765Sa+yukHqz0PPglCybWhmvXffBUy4tdMoaH+G91Ofc3l58ZUGy9DLGFeJChJEQ1T
5WSkY8LWqVa5vGl/wovBeSMVksXb2WsFPPDpgy6bSX3zej1PIJdOMWh/l8VFj31rLiFlQao73rx7
EuRtp+7lDgTXjwxWzfgFwmv/ht+IF7bzqPWclE2IsuPFaEUlgZ8YBTF53u/LLPn/VOZFtzQKGqDV
Y11EJUNJUdq6Q57YDvSorLICca7f7YtJKBmVJY1TE1RUaZ8FIN31kH/9M/w9wlVUkL+U/EtgVGgo
lRBCTlEUV81udgpt1ZfybgjTs+6I8iPI5GtyNQajuFuse5pLFnbmSTiuizwKJmQwegAvLJTNWGry
owABayJ1dEYTKxDIIBU0iYJQ8HrsQZgs3Az9P1nh5cIMbNo7tjn4GFBLaUQlvaNRQUeVcEYM50kK
oMznX5ZraPmDcI873ipfPmiadfBE14gfW3diZTE83FteUH6EYf/6aKo+WMaMJ4iu4+4ZFcUGWIZv
YcyeWayre179EeIc7MgBCa4xdBdx5ty2eQQDqrRVns2ygcU1siGvgYy28PWMfHeIFmcUcT4+Ig0j
9Onn0+sbbu3Tvzoz+xf3E8dif8arMJ4h4PMr6UcRAl+l7e4xvki+Aer00mnbBxchfZhkE/OY/cYd
Wjql6x+l7KJN9mFwnLi3b8uQcpILMNLGQ9AAeKMIeQj2BQFb3YD1DsSqe9i2s7qqUumoifsGOFXD
yf2R9f8UC+qC5yNaIXHZplcrJa0+GyqCizkfRx+KMv0BUQ5Qf6W0EivxoICc2VcgJQBFe9rlKaug
FzU4bY8s4QMNFQ3/HhbSkupccF4ZFpbRkxqHvSruNx6013yBrySUQWhH0IBc/BmLof0V4k1JT81k
Ql5uWb5OEGf8PLG84u+GmPjxJTjH/0UImDAfypssmQU19nQgb6vAZ4xxhycHZcO8Zrj1LyEMAgah
T4RvlebAH34JS1qtpCzGsZlFJq+7z7NSR7NNnOSrwfL5RnfbbzxcN1fhrwn92wecFMvVDOo7RmR6
4o1sBk1dmLANnbP1zK8XDZSFQjAzWf161b2Pk5iuO6YwbeIt77OLlP0zhgND+nbec4E4qCcGpg0z
/AmLw3r/vP5jA7exlJQa2pKCHTQgeW5CWgUZC9M1gQTHp3eCnMiJUnVsILQT7nOcSAUXKnkAW0UI
50LSjpI5bjjuxZHFVG66oMWEOGOyCvHXOi5cpfUtpIkrzVuBoeYyPIELVel9GNsUqiUrsLwBZH98
Cvkddemm2Dbf9ppGH8tUm1oP2tn42tl7wRluYWsJF8vP3vTtGpiNRhjpm0PqdksxzmWXbTAc6FXS
bE7sbCvAVE7OZJHyYfHVTSae7U+nZ33Fgrb4Wsisvy8qxloXKgDEgXUb+qJCHFDUjQXuZNIeVyaw
iEcX9YiBIaYwVauJbp0EP6a0AoWxROyeTBvnAILJBlXk5e8wePaQqSs9DCDdcjrHY3Q3KRBJiFE7
J1Q+OdhHeIhlLTuFDWj3Z+ejaOwf+Oeenu/ZRfK6AamOPzWTkLLEsRXPKLU0WmvadmfPWEJ+BLxk
uObX0k4j/o2CpwjJ0nDjm4Cwbf4bMIE8a4b+pXxKXmE4KMYL2fjiQyh3zzqrm1pNf49mQayl9r+K
Wimu9dWPRWQMJ2KW/nuFi31vbUPH/mJKPmp9HWDBZ2HhEXFFTb1rwBgLLFQfo/xwhGfzLAw1PZp+
NPknI19WRcl0Llbrldw0BrJSB0nMIS8T8JVC2KnkicldsfzjfAuBdelb+cl01avTEZDdeIXF0Kap
dihZ/Xotm7xyvWkO1kyN/W0cVxWmnqaXJZ0nW6j2jS2KZyqE7C0y67AalDG+GabCwffA3c/gBbQC
iOi7Yw5QL+5XVYU+V9FjNyXU3EtCcrOvEpFMbG8ikJ7OX6YENDsZubj17dchcV98wbU1YHjfes+X
P9HvRAB3b7j6T9qL+YxhaMnIJPWONpo/oypzXT7ymxUtzdjtl33AQl5FAgsQM4vwKu/NED6W11Yt
pi8rCrCk15yTmaXWSJWJgbVXOSGFFfhbSS0v5vw1qhSDNefEZNzmUXTjtHf0IhHsXs1F3jgHVRet
Cpo20X8KlhfokjUbFd3c5QRfjrJDfHhQOh9plLuBaOp+hZPRY/m3R9vlKE/DaZdcnUVwYuKAyXb0
jbxJcHbTbHrvimlQQ+jQdM1Jo7jimRHQwgbU9Pofwo7hK74jAJaf0dR70xZ4q41Ii2eolTKukdM8
g0a9D7M90VcmHqZ+3kQVJNSGmvJ8p8ud/D1/Ri8ea9eIa2Cb+Px3NxaU1uEjkYeRvAXRXInz95xs
4MLf18J4sMkFuWBQBGDXrEbW2rbo3M0VjlBOQtz/IipTZwn12t5L7EWjTZ2ZzGX2H8sTYbuX1iqp
9KJxUrug9VhBytQdsUKXqfI5P6lhgmzY12OCPx+I9jct034bVo6GdfaOySvx5i4MFKAYRI9gmB/M
R7l7FG1+VUx4GztTXZ+3ZX/assWE6oYRzm5fNwHVABy7tCfn3V1Jie4brkODiS7t2rpfUqBelpMA
czfNu8R6sIpadpFvQa1SeKxhvi2ogRZchvp61d7cz1rK9Uk1mdmMVJsfY7z6p38x2xN/h8dLJvGl
ViiGtqTw5URwplehvAizm1rUxjWPAHYyswEUU3WVSVq29TGm3i1JuXTXMwYdJsJBAjLrsmT2uDu0
qHmX5LuWkFkM+SwmDpU2Duqo+G8wyb9RfYqh/Hcz41nI7q714a3s+Hi5L/4iQb6OX0Z6PIGfmKid
yIf5epHaaz/t/341a8lfdw8SadVm0ZJihZEp8c1Z4+NiSJLCbzKtbBy/c1k2XibGwhdrK0takZdG
L2ps9SfpQq9fNgBedgCZcyHa85t4i9lfD4/GhkrbcQUVw5u5pX6Ffb1v5nj5J+TctetncN0aKzCb
Ah5egu8ogUEYIwZdK+o7rvyufBy5KoziTUHcFwsrVQ5OPIAFr19KeBje/HD/s2xl8DV/P+haQNja
utGh+zQy55SzFcSM+Qk3GVPqzAmhMAFt3Zn7PKdl+TwsyJYrHdbODz6el0d3VYblf8dhjPOvovZX
9nnACWjRAoTzsGAal1yJTXJoAm0/f+oeTSlgCsm1P4cadLwpzcFYNZwpegwYAl0I/aJh8/eWAu1s
0jwrJCs+YKmW979RwDVfG2EVLCKCtT3V4zEWp6hJTAY331qYXpXoIe83VrFmk+pSbm3GUvF+qIb9
++VXhXjawiHeuGM5qKOjqRZQ8tILOZR4BT0masTwcwEwLQTSVEzgFe7l6yq993rDEa/RB+dHYYwf
4psQ7Yj6qxvUKGtPAqmQJIXZRo6sU22rvN+WrTDyTQsSpEPB7qwndpbYlrlvmGSXiOWLodlmHgv1
n1idyuo+Xi6cZJSF2DXbXVHY6nSKtvcU5OWlGbqCIuz0AcPSA79+2ghjm3x9CbfUE9UWvIFfdgHX
qyS8RuspVH0SqW/fksicBNQw0OGfuXRMI+36C+4oVyxCpGpNoXqBlvc4suqYbR0UecUzbWkkHZb2
602a0oOSrpr+I0gQU48VkHTw3ILD/kiXQk18m1CBiE6/YlpxeEj9v6SxgZOijcVNOfE/QY88jfSJ
UeacnmAERkEr1F3bis8owG5plXJUmIoBRSDMISz0lEds/ch0YGeUirwVs1Wv8Fx8j7jTPg3LWTeR
5aN3wF0yq5tHMjGvAa591jl+joLFupue21KC808iJeBrVPxcY593cP+8TVGQ/SrDETPJrMwF4tBp
KfK9aM599LfifA3ZTp9fTjX0CsqxHQM6CUC/e5rCJ/6lTVIGPTBHhQYjB82OnzMWgDZTI5XcDeEz
7UNHwcdYfwwsOpPIuN+T4WCFnzJl8o3FPiWGqo0KF7qML0ScADe8ZbbJPupFaME7yoBU4EznPV41
FR4wllmLhb9Xncr6asaGwvBjQ3Oe7vo3Oqt7vhJVwYMqbdtHLN2d31Q56OrSk0JmJfpOZbQ7ZbWz
nqZg8fUVTkcFgNKvd/emgyhirxwOoS/SJ/eY0X4Hnif0Ofq2Il4i/gfTo9zA8/VsaeWORCsYyDbh
XxvCGVa/ZQTxLYrD5Z5mEqxp0cG0YMt48zlpu2SCiL68FG49/YwAi6TanTsmgv+OdQJBDXSV9ZPH
eq7Tm30ZzzUAkRuMe1BBTk7q/APbP3eSsAxdmpmIEAqchH0wdGvS1bHwgscfL4lGC/cCki6Yd/sp
Bws/szmO+9l895QF/XPcLqTJaqaYSxM1br5zlLuTlMlFzpWLSqWIGS8TTPB29Omg77OtwdJqLiiW
3U1f4lDfBWj0QSDzL0nqSCAA1v16X7iFX9fq8iuN1GMNPJ5gVOnYzd6R7NOj7pz51YwyXPo2f85f
FVTKE1oV2wd7qzZFMUHG90KYwuDTw7BRRRrYwPWU8rypLJ2S+H43g7gJyqu3MAoB9tsdw6lviCUd
tW9H6s7g3u+2heQSJFgxRquz2d0CiKKO9t2hYF71pxONwDNmTGxlqTCgV4dVOTXTZfEcr6pvpRL+
1cHJqjfRznh1l9Uj2J39+XEZSCGWxrqNMLEOiqsNZnaDcY/MJfRS7Ar5o6hDHwM7/nykgU8C9m3o
CfykyzWqD3auDBaTPkdh5rZ+fjfBMQmEIsYA1Go8aFLjXJ/Gvc9HGlkU4QXmQGr2dXOsXRdqZwyr
dMgpVpOVT9EdOf3mDIbm3KwxNyzkxu7iJ389rKzgnWoJogzmDB1oK8kWVwK2IoaDP67Hc+YcR2X8
auQIPBamVXCfwy7TFbYkWUJLfaIZSUhpO0bBc0qWAwxtKEgcVR1++G3fMwaJ1uzUgPGOSZuRmSyu
kMOSl4/KekIqbgixRf/J76YLVjgTMR3H32PWPtwAunRcwHKAhL1EC/wzQY2imdtbz8Vb2fHU9Ozr
2wfuuhZ2HS4tRZMEh5tq4765GrRT0uSTvyOWi/JCO8g/5v1CDvnTWtDgpqnyyf4yKhjAtNMBXRR/
1Z5T8ZtDPNNnH2gUWlCmi1YQITcjqNWrHLUgE+MZACQ76veb4fW0Y88QUZ+dDRRMa7ThEjKxthPO
IwUraCvr717tzzT6iP6fF5F4G4dnXLto6YF3UwfobbTL5yZiWXJ69jcrdW3iO4KCzIewvZ+NGep8
ktlSE5mthHttAP4rRoLR/RK4UCSz2L+jh9iEnWLgapQxXkoChCLypHZoxUODnTieN6o4PjNA4nkT
+EySfX+Tnp1zNm5qvDhRMYxlH5weuIcpouOBiqJHAhFxiszAZj8GnyABmIPx9qsX+b1CyBwVdJEn
a3YIVG70dyBfS3UjqoWdSWfLVBESFKOCHC2a9H9DG2Sf/fFQFHMSN81lJzwwV6xNoUcluFA5nquF
G7AP4AvVvjdqs3a77p1fP2RphElvm0VYECyBPNpcZt5nFS55pKYLvb7G+OoreWnN9qApxbczRYts
///6Za4CZKggXvZIr76MOGOI95V3x/vlKhZjdDHdljHZECCziU54T3RlDLdv0bS94idSBNAWmcNL
DncpKsYzSWr6xytTxPC3RwRT3tiqMttajZNYvsD36HZ600vlhnIvOiNctV9h0OHvzCWB1GDMdnb4
WqjVxc+YJLzq+Pvcn7IKAfGe2Nol0ZzBnopRSTeBTZnP/tb4OW0v3AkEsTJT5PT/NoYkIKEFrqWJ
/b1SfGw9Nb2i8Bh4unQwAndyX2uGN2ApF5k4lBuxfEMNUrlIWWc7omGpuE58Uz62xP2oo4eveu8l
bALpD4CLGopECKq2XrFke2Ccg0lmeGP0SmlG/BdI6hBIA++hsyEzIq2WFVY5+YBJj+7tdOBv5JM4
Z/iRKMnvuapBn96pfwgKqDrRvlVuvALMQ16IRFRKOdBK3B72sOh4KzZi4yvBy7TQPBxgXOTp9x11
rYC7vm1HgZ1PDJZ4uOSzNBIHWhTv3zRU4ZF3Acay1HFE90985U7umZNDYKa3MaG92nnJIPzTFbtL
IYxTvjfoGF9c2+dhh4laKaNyBMwPOFzu/HdSyLRprI4SFCLrPmllYeAhuGg/fsdLyYmVTh2+9QbB
HH8cGHyJdR0X5hGOMyyJ2cHNc8cSKcbEB5Sf9SJp2vHY1xl98t7sE2sIFrGhr8pFeL0SSCqNTZmK
PkdtV9zgkp4xzw4JEsF6p3ji6u+DfL7w2AWcHyQV1p1dqNzSt+wHGOyvMAAxVeSFgkjghGdhThM/
y3VYM60kX1L0N4jMF3zMdXTHtwZkBu1VL66YEtBzod86qeTYGXdUkCSqXfEjUJSw93gtzSiUMvwh
kMzZ3APr6T0YB5+OmBoeci/vLWcQ25KBDmHB6q6y5S1GYSZw/CKQb915P5cmqlRmbsCyJOtIr+nY
jHtrDcFFrezNmVj59BK3ZRwK6vvlFZMRrZpD8AxvHJ4mTqFvTUhlgaVJ46w7fq/fav5kRHFbEEfv
fzJ821BfLSdUkoiFEY/Ik4tQEB3oAdOBqs6/74ePzvOIp0xAitfW7hEz+B0Txy6uipgDnzDI9pQa
rQGoa6/Phh6DxLN9m/MGIJXjo9BSD6qg3CvecuN6FluUemrzenu0qVArQrLwp6rOlbSZA0r130f8
P6SiBfQqyAV+N59ZqGJfJmp6CZWt5t5uhA932VGSHXHVQUWlmiSnpm/7EXHF+R/6EeyIT/A8KF1g
K/VtlO4GiM91PehxF00bG5aD3ps8yDcla66LNM/DXWpWKrZ6RZSXRgu8L9mWn1VkOPCssGool5fi
SH8lIr9VqRauJwIwjwSXs34BULE6FAOvmQTxUOWHkeyr3KmYRmbQva06giOgztwN6hTLP3iMTBTz
YBJVWmOuXFaSe1VXNlD0rbWV1xjYHAcf4VGGSLOk4EKk5aT9OJMjTeqrHenWnbsK9g1UUaL+l7Wi
sy/qx3yk5IZkJvBd3dk2rszCnztgU2bsjxvuUdVuGTjB4jSEJGlMVsjxPV7pJ+6Mi2oDtsAU4Unm
Hn9p0VJd7ze0QgGpTrcQNn4cJzLGf6kI3Q/zlIx0fE7RaQJSdlDmWDSWM6ep5f1+8fsPfvpnWPa2
jWzCqORDsomglQSynPXV3YQxVGaxoT++pCQauyGNzqgUz/2NZHgxu1rj/EhwUIDIwxVw4PtgLqzx
aOVVI0S1g+mcY2y3JOzuGIqKi/as8nu6/xRVspY3kpxi3ytGGtJ+fXa/jJPgYszml/qLHqswFDsc
+TbxUhEvhCFmg3e7kwX46b7uA2VVlc8i5mVPiXIkcC3J/P3Qt76lpSGufPZFE3N/wDVAb+hK5jEi
6sgsrLyFUTmXSyJ6rbKE4YjpZG3dSMZQ6bWQdXwj4wMF62Lby5BGV46Do3WYln1gABsJBYq7qzNO
kG1kYNpaPuRgh4cHgVnW9hfVvO7JImj1/Kw8Kqh4a69WZuNfyp7h76FGXI8NIaZKPwF0zrXkE/nJ
nNZla1wsYRaT/rY/9cM8ZH6Mk6IoH0WyL0nTwFL3b0O0+ML3s+nl0S8H0h7N817HyDQ2myqtmtbS
nwoD/WrEMZ/k3LNHBZYnOgGSuHmWy/0lTfL4IjmdBwhPSlBGcO4riKZa75I/oIyWEjVkRKMG503h
+/AoUraPw/eBR9Ep3816YXLr4CoKEG6E1Ei+Fd4fPkJ/sQGNYPc6gL7LulwVBU48/23ZdrKfYxoW
id7sfweHFRvVS4n34iwHj2IFMtCcGBBLUS8HYUBSV3vNgNpPDL3plRWBwpI+eh6IV6QCSUttweDP
yP8jH6+VPqPCNoGx3nqxoz5MfEfK07E8BY/zKfIrzam2y69rbVJ9M3br1HMe/XGyvc+SWcVzmMcE
yPNGD8SviWPhLdP0m2vGBADh9WXsbboHzOEfh+Lzzm1wiZNs19dpKvKRCV8J/SBhldP/AJn96rjV
j/j3rqyAj9okFp1fXIEVwki3xai4MiJb8wlpsdrzRPmV2Q/yFpWKSlEMJlqBHEe1JHd/ZS1JKR0u
bInK/msQC7MageSufJdU2NkjwSSslVsT9fm8EpqiGwmSZnCsl8UiNlrDYyUHCsp4LXeUE3l6hyil
mlENiEsxG7AQNYg9Ri1229FpRIFDpECNQieq039c/9wck6S6K0zLkNkVGWQvc0UyTfyM2NbIrUIn
HCnHeYCe3JoWgzdzhA7ZFqi8ZzrIJ3EPkC7CHEQPgQbjODfj9ITOKFnirQGhP2ehLvmd8zB55rIy
pvEF4OO9ixa+B/v7N4eqIF408Bjmi92eQ397pgnY8s+ZiDkvGYU6+0qTMM9kDE+e84f+gdId4KlS
YsTf51jql2fZBu9RrcYhsZD81RXwUfIgqjTaSxx7x3uuKvSxL5X/1gz0YyzUCiR2uDRWS36k79P1
bTGdl1oc0/xZrGS/vW4ktgHfF9LuHiRTIMAC/nA2t+sqCZLoVbtlDBXFi4683Th1Ym2zvKd4aWlv
58zQYM5m50tE/eD4jCNgVnPB1VTe1cTL7rjIFMvG0tMQyBibG3lTSImrn1SZpdXKRKavp/SgL0yx
FI+ldm1Aaa8Yj5GcIoj6aE3sil7q5tu/oGORD4kE6RxqSPJGW7LpVBHG8F2IxE3loPuzan1LV81T
NR9A7iZNyDtGLbmEy0drvvUwmHuo9bMUKZZZEGP2tNtYrSO02dne4LUkwrgsHWDan1xi3YU0eQ3P
gXyxhM4HRqFMLn2apcpbh9rciBnfeJJaX7NR81TtScTTlwOQNtQsv/Skm0IoGE5zIya1FJ3Nr42X
ATg7Z1awldU4wo02WymYTIR6S2NvpCTddRYvOuK1uScvdYpc3ooj/aECzQWSnTiRxosQX2cUex+U
Fv55bOcediXzykrHnh93ahnPm+MAWoMT92hNQ9ipcKVC+AzCSXnv8MYt/SDN9T6ixS0C2rGNmPdL
Y4EmL+1Lkv2RR4jgBRKUjlgurO0a8d7YF+BP+2qw1Hu6BvI+97RwPF+iotxB+qIlKRUIEMHrmMcy
V5OIjdnTzhLpyIcXycSRK9Kz2ndOPb0r6BL7I/MHNG7UHwk9aypMy7rWV2uw/a64tVAh4K742ppj
jyc86gLnOd4Ibyg1bPajTs95TjGCP5B4M/LnNsGejX8jj7aHu4hoDKsKFK0sC+QDDlvsD1ckJVhI
uAxNX3qy45EmB1KHhQ0l8yoOyU9Rkc7mm44njvKTaU+VC9uo9P6FzS5QZIzjrWumpP/RXuUA3v/3
9gfSBFMMYZ6oJTsRgvHTe6bGnQhM/TUBzkIJXh4spqmDZdx+Ih5ltumRisrWKMop/Gz0/ptfJWhY
cMstqabTvi4sS5dGDcherVMGoy6W/uo4YUbv++NSB/dT/6bNOKRAg0oDs/Tnu4T59xFOcYRCRrY+
k3/VP8jjE3Oy7vUhsCzQnQJKzg7gffLyUFnzFY8icUpGjDIcDxACoa6Ivd79+HVvEiGrsRaAYgkh
xcTA64WnXER4bgEgvoMQs89YEf/mZ3WbWPjOArS4xyUcxt3weUohXel4GsZz/+JdyaWUR3k0oR0W
a7Vh8LLfbbSnQfDauAaLQ1hTNziPh1XEJj8ZcNyLZxHGQE3dZWLjwFVe9cUNMxnMgqQntL8V/cE3
c4vA9ABDaBvQ7bPvh6fJSp+9SHJYDt5DAWXxI+DJnkzVnGcEQ9M6cdt3bX+livaTSAQ4p/0wjRqR
cEZ96NpHGwu2RZ0RMJ8N5LqpZ1+Ti+lncq/bDCdhud8ENWJz2gfx+L36Nhi3kubTC3cwV0oTMYIa
TmKY0Fi+srzp4eWsKJgzghTYipHquzMkJGkk3cC6RDDFoJtGZAK8AOLBrnsWvZN8sjjIDuW0Ns9/
k0iNKUYQkEwhWdy7d7OjX9/GAcnoovhNuHAsJ08eduPvZTxT91/gGCQth+TmMrpj9DM4/zJFAX+Y
bXxzRZcl0YEVuqy3S65uAlWgGa38/y8wyHSSQkOoNXZX+LrEjyS9mUzJG/QH5+NEzpEdaffZvumz
Qdd1cQ8Dt7D37srfEOGHocV7DUDU4pzLJ2NCXW7b922Iq9K1Tze7doWG73WOmVdiHQnfOhbQaZFP
5Iz+fXFEHWMwzK+HalaEgoPo6TvXpe8FmPR1q48ZeFJM43gaEPemFyZqftXyhV8iRKnFUvvpoXgL
L1gm0YZrEiviqMtqoAhnmbR/pPNuhHsSIuHYrSt2TTXXAb08IOoJDL6uHXfpUO1njeXsrGKD1SrO
/ZqYok84TxhO767MrWKCG0wa9oX0G6JMKEjDzmCv4gEBEAZZxvV3BmKjlOxHmUc41G5+7JtkTrAc
JpiAKRrck7Bj15Lvd0x3+vffjnrlJ3WR/ns7fFVUcxAxwA7y+p2oBaV2TUbr9hj+458fQu508mrq
Fa7YoE9vg1e+HKEai3MSDIAZdZscbcFVOytdwguQ6Vx0IpwwA40lbd6+bNCAKm7CA9SSttFjzjXs
ssupd2JpNjyBTEt+rArLK9BrbwIHA6O+VhBI15WCOVaNvKtAa7aNdqQO+gg5JHBU4kBgseZFj6Rr
RYHTAyWw0EGRF4dkvpPD5PD7uN1/mFukR3F0+nk9VpaTfCG98QLxvTiDUPjguDc+OP9/MGwoxvT1
9Z7td/JNTA++Ugl/lDymYMRpmRxtE89COOw4RlXNc1KRmlFEn4/qmnwaFzPBOy8eWX8EbeiKCVrU
K8T5Jf95shbsCYk3lqj7Q5hY5OOYJYcNWqbrS/yKMxxa/zPP0TA/PoE7oHh6yu3mZvGDNlfL2MSF
h587mSz6R0bPEmafOxWoT0H0PlMQ3s3uLs7IkWMkJa0mAyVq+WXF928mcr1p16dP90E2hOw0+oMe
e1XriCWArIrcdAu0oz2La99QDQmL5Ir0ps+nVyh3jXuQ9OwuechiFitSYx5MJqKkgeyJSRUizLyQ
2sgCDyZlZDIr9UHQRFJRQjgvX2DHiSKgC+qt/OoEsv+hDznlNoZXSjTeqhzYaNBdB31knjGXfke1
OfQ1u3rjWN6ksWd5oSX0jYCOprP1G27qSiPIJFKOfS2lltxpy21ARuL/qcm4uV2PB7aMiW2rtBSO
ok8dDKDtube8hupfb7YuAXeAy2MDli1dAz1oc3iAQ+2G3l4Zr7KWWHyCy3mPPf9Jy7aaBkK+WR5v
5KrTQLWQL9zZR/hSXySu64BS0Fmleao3BBCqchIhYV1rpMKvBuQ/sY6AZEyxxmlaWcDMsN5jr14z
tGHHXuIJ45NBG5zAcZqSrPGeofCiO7l7iaA/xFq9HHHaQuwij9X+vfDQAGZ+MzHFgQpEBhZWjyCV
ow5eusJDNkCWA1/bp3J3KAOMFPmsptQu+oz8s/8cZGvJc7NpHY2HyEnN49BC4sY64YQTz6z9hZ1F
gYXQMOoN9mv62fjH1Uuo3q1Cprukl9GSYvS6x26+bCa/X8/31wPR1Q7JorWs6hTRxTcpEQOLOEKK
9Hw5VNz5xMHB9/OjdZceFh10170Qm4ujH3fu2fiG8a+GqIJHqe20qXqCN4WL8dijfY50jMIKD5PA
OL5MgQEdgbLq/iGr3+uWBGkCU9FgDf7Jge6NYWMZXcBDYhR6c4Kg7aim5bcmnFICF5qC9X+MsbeM
EEGyFLd2LuC7HAgizz25OJTTIYkJVg809HQQ4shewrAQZ/G4wN5LyKXEt6KIMsU27ddHGD2xjtuE
rUmo3tBV66B9DH+WoBVNVrZMcRt3FVOa7ibG+nBI2vDY+n17JQ9ICL6nyzmKg6HhCtSdWshJgwiN
ESmPIU9TeE/ybOBu8X1RoGIPuh95iPH+xiUl+5PdLX9gVQEcmKp+UvbYbtlCfpzcEjhvxyNDNNtS
7PmOYeY31EKj0CK13alifvQmbxV60pwByByzVRbAfc1Rkm43RVBCfCQjvGyQnXdEbvFzaWRDrvlS
lNneDj9CX4Z+L5JWBqJ2gis6bsdPppruGqNBml7sO6wM675FQV2949YQN2P4/CTUkI/SEdw6W4pN
vHW+xxf214m6I3+c3986n/SDQLUtOZhZ290R1veO8sQlf26vbODL8bpl1Ed93zdNdaL2lKP8RVbu
EDLzTyuaXGgjZ7BJIES7F4JaapjTnd7P8cJQyueLi/ILrTUlwF8MW5hY+StOQX28oppIM2fL1sct
DXH3NRP2RAK2Khe2GQPEEl0t5rDYp6ACqOLkBsrHHt9zg35Pbzs9AvBnqZk9kKZIaWLkSTleqcbp
vw+cb8i2eC/yewnSJZ9SwQ4yinvNem8MUPwfVCfJW6IFqI15onhQrAEDIYMeDjHkMk68KKcf1loT
YJ3Ocssi3yjVzHzzr7JscXqcyeB9IV60G+kfzDAnFN6r3ECL7bDqqxAq7/umAHCC6HIcKHHp1t9s
RjtGDza35OFEq30bKm6kK8mbz4MEJr6PpEffF1+KhVHRM2SwvbBBHBDZjPM4FaEqtOvD4SoX+WMa
Q+eQMWHZa/2gHV4v3252cg0hrwvGwngWodtG3MbqGfou69BsBDj22db98ZuxZeWqd522fQoF703H
oRricMXj7UrWOa206m+32wZf4XTUSnek/TwitA==
`protect end_protected
