-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
W56jPwMqvs3E1sInnH4+4C8/ZrJUi1vcCYBBvU0eRLvImRsgkqd3ZB+3CN9kbF1Zq7ubDvxaWceV
Yql6uyVmfZNMygoKA2O6kApAZsQ5Dm7x47uma1m67Kbfa5AEVNAWyNZyvy2ExUnXoBC+lERGxfRC
QJtGPLaVnkl+V00bhXvOrEKptojgUVhOAYU0oHX3ewr/juqrvI+YU4T9O8YzHdTFUQaeE4FjDU4B
Qyw8LaecxBwrHNInbNWTrftFo7Dgs854//oFqz9EVDiMELH3xF031LrWHNUq/MU4GNu6rcA3mkW4
YlmKpo8+Euaa/b+XvGlxgZdr8n3pIeerwg7N2A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4448)
`protect data_block
aub+cZCJsTSAXp3ULGV3hA4AphTGfyzlLMoOaYyWvb++RA1gQfgaKm404LacsrLydP9wEYghvebI
k9YXQUoS/AhdrbD69PV/LGp0rL76Q8YPImbfpAhIK7tagJ7fE8kZE0iVprB9EgYVx7CQJl+V7OtO
bis/menQZkLoeqiAxrOgHTWslrD1BQmQtrPlgwk4uRDkBSODlcf6HCPXSR/mZxqiOvUcdtJOQ2Oh
zSQDBdP8H14ACDT1KpgH2otqp0Lrw+8QJk7FGI5SeL+I30i8fy2rIW76MUTXb4IMJZVUY3VSUAid
yZY5WXQv77f9/ebkKFNAshKcIiNqH9o1ENBKxp7+eNqLs4ob3B+Aql7S8OoV5yXls12xrjshS9gi
qKtho3xt/ftsW8DJIwmSL3YwxicuWwpO3hhgy5V+eA2oz1DJk7NocYP/c/LyZB4NgUOCJRRElQcm
cmnf6k2HVmd9OdDFJ8F5P/5bQseDaS5Nw+0SfuGP/RS4WX3m2Bcj1WDDlGl1FrICE9QsTULyHdNx
Uwtnh4c5o0gEjG/cvb9F/ByhUWpUFQ5fRxONQ6w2xq8Tfh6cruo6sI7ucT1rWHtgca7gGwSVUaRh
pF0ZTq36tT4fKMULwcIUvKZJ5l7nUn9nx4eNzf5sUxexv7jdwe4WWXXifOB/AW8EKVqfC/AHlpQH
iVKY5GSRZ2OK3tQdMzaaocIPrxNtHRQUZ3driMeltxIE3JgZsL+MCxjz7uzON74AEEs6WFAbt9ON
VbrWl6Ym9QIYJtPgcubgzVoEh7c14PEGuBfDR/O5sY4Ik5lRhWxoYWvPaa4aO3E1xK+o8vVJh868
25aGK6dfrLb0nB0pqlDrR9t+Owc3nRu5BWph9Jj+kKQmWn+PmSowOonZxXB58TRKaFivWss95lo1
ynDeUHEhkUuLE7NJZ4JldE0k6mICM0hgPAlO24hhnNWsNjw22EIXDSO8PKrNHmFaEUDrqbMCM0d3
YbUswEXAU4QuhKP6MW2fnUNFe0kwimNECrzBo8MocBPyTth8ANqxBf0lqQ2zv+qV+1MoYIZU+Xy0
Kpd8mAB64z4WknDPxaq3uDX8Ai9B8AqbioAdKUTxjMR/pqHXRMqkRM+0LdnfkDuNqzsC86BQEZbX
02E91mtRd+zqrEPZHzHUK5UrFu5Pz565gfmqFU0HVxl8BtyLc7xZPHaDHlWq+kPFGtqnrXfBbHD9
VpmBOFGik10FxivURpOuTNaZZOinEhZMo6rd2/BpphhDSYxIKyZxtHhpwqQzPA6euf/iXbV2qpYC
74pj32OX9Thro8LuHvcNSL2JGb6S/c5rXxEXaLFo+vP6kD1OR8rj+dZykeZrK6IKAS4t5KnlUiIA
dNW+f5MLLf79n2PTmyrzP/f0q+/avHvXT9fmoc/207YYoLoAbYTavqOtyJqa42aOl1ISA1GcooH4
AJTLmV3DGYnTJvEA+9c0yOfj0CW9gZMhsr0kT4fLJFNf3AxV5vy4nVia3vYm4uJqd0osdlKIau09
Ok0615KzddzaOwryitSdT1mpr0IoKYJXkgp1v/EBKkDrf7Ykdz2utbv7Fst4935H2hZxMfk3NhLX
9dpVxrRaxIwsg0hCT+kuXnUYr2tN4TjL7D+g+jfBW2kc1fYmzp9ke5+a9vHmaCmGgR/6eennKXNv
KiJZdVpfDTt3jhykAJ++poP9vgazl1HcGP2CUr8GTqgaEADj5H2SesgMqH222yzHLeOrP0mEqTWb
IUEBzlG0B1BFnkchwrBtZKdIdPOTQjU5bJ/x/D4cFY8WVb4xC/LFP5HJNhIRZR7Pjlt+p4YolU1b
malPfCLIrh8Se5vSZxe6HcIaUHoo2dX2lmwYi5YsWdUHcx/wXPUmxcVjSHAyerYo1a6tsvwh0+jW
O3cqaoeRUH1Fyarsmv9xCg0EKpra5z4i03ijC4FwhFKpV1oWBrEUEaC3ZogoDYmyM2trwOe96o5n
+SOAnvVG4ZF2zoAPnilEvXkshNFMLjyx5GtrICAX5b5gxudf581fv58SxoM1Eb3fg/iMuVeBD7mA
Jf7tex+tNw9Pg50Z3tVsSKS6YASd3QumS1egyEcdh9ag9trK8UX94pSMINEWMHpE0XQ64Ph6eS0/
ZSwgqvpc5ik76d+jAIPPZjJzK1aa4WvKyra8siS9MBdP/aziANopSkxefEOLXJJJlCw+tvfiT8CJ
UKtK3wFLwMMisqSuWoknW//J1prWVZcMFyFa8EWv/JCqXAZs45PyQYlf6ipU75uZWLolck5X5D+8
bwZyOxT0BAMTWUT2t3mn4NGyDrM+MMMZb9YKfoc88MssAN8c+pdKXeCaOn6voa01hmHXeNXji6ga
H4Q4bfBciFpliGUjepcnqVwR1K2eALIewsKaIgC0ITEGjXv3/jx58CONyfeMKglOAdzy/WNtngsz
gx/3eSK8bU2JE3i2pG0Z80ru0OMU8X6rvCIqt6xuPCFbfLvefTFBjUuhwO7G2x6xDYwJAJkFjzd2
ptkfHKizNIh9AnwrGobEcbtadgi65PSxFSLD+NOSmAl1i7/lHN8QvbljZJojTzEkP4INbXHyV+Hk
S+VcXeQyvSCixfA2pn+Huo1YaA1/Is+M23JGEQbjKYujuJqUpSHTnZqn8PxO9xoSRDQ6WzG4d7ss
gCLj6lCfzxy+wmwqPYjCOSCNI9n5JqaySbupfl1uJOQXQDOpohQxdxz6xEF3TMYGf7a/4Xmvj3Gz
fucFNiJ1CQKpZYNzmM532MoAm+ncVARxEkwVYffT+pqMsRnknhul+PCGb9NxzDGcNpbwRoWHasWP
+2paNZErN9Hi39HlYvXrDCooPx4xKMxjnUChDt8D2PErvcb8wvclqWFyRmCFTZCaWJUk36gaBOvv
xO55A9ZR6JN2s6wXpN3yT+uUdot4V8I7n+ME4Yih8VVdHoaNYdUMDd7CZSdrzhHf1+BF+fE+CMhI
UstTOl5aLfBRizBxoJF8WNxT4uX61Va8bVEESjOanb/a2+svJbYGkiN7pCQsXxEYlS3XOWwyCBta
sQ8GmsGvoHmxpzNtHhoCSJb9ckcsDT3BHKsPE4O2YOU7fRlheqh8p7kq9koYRpgC7waMXlFTHj3c
1McE9uG7CR229fvxaNqxXc2Hw/XkP7KM1+DfwhAMPGYMa2RTyb3PaZcZMBIpHSD2gPNMY3X4Zrkg
OCweSQP+yBGWUyOGscFpYzPjINDB7sAarU4U6b3FllUW/HG7gSNa5IpTiEv5lmQ+jYxbc5f3iE/t
HUxyFHQ4kgYFyg/ZjqWO6YDKK2UahkplD1JkxEyqfIw7V3pazwIzvdW0nQw0UNEh/6opmPBIWEwi
0EOLLcbpwkwoTPWvyp280uTkNDYnJtU1lKZHi5eUgxIrRj29wfySge3oQ6ZMD74t7eEYY5BcRGPL
WIH0bdkGDgWH4fpOoOZIG1F5b95FNh2NqFth1Vo6fvYCQPqfjN9DsN5mPwAT/O+SSum0V8jdw6uO
hvDM9N+J16epqD3myOUtN/sbWMEw1Q//8xbklkh6iwGXALK4x2MotpqV6hemcuif5XoJzSHX+RKl
5yMXRpTQwuNl0upDgJUIGjgweou6RkVTMvzXwJZLjEgMu2m3AKCO7VAswhymwrCxgbVzRKIi18Dw
gawQ25qKYF3PTXhSfFu+KIVDh1V8KIQ7+hO1gqwAZNmlLHoXp6oYivzs6uC2noPsgcyqkphT7EwT
B+H9qJ3cMUQigRWGUqCNqENaUDRVf6Bw4i9iuryc5fVN7QQfKtZLScjoCqHU34Nh2LT34iwkt6sQ
cLE//Ar2zYttC+c0ITAe2fRPThY5YuHBfuCF9F8aZZURm54xLxcIuQUxOW8BK4jCCh7DPgHlyWiZ
YfpMSwkKzbhIUflUWckShddVEE/fR2DyhW2xbDBWVsnnserbwTSvd3RWhJaNqfReNhww5uz33rxh
doIeMVmMj6kHoU3lMVC3QXC0Rhq8KgqRSeLWOtFdEdHxTYG2n6DNqQ3rO1K+pQCnFfyOFja4ruk9
/8HrDlNqYvzmIyRgMTgUiprxdxb1h0K8alcUXh+SOZDMi1/pWyVJsNTCpSXZLd41ztOgw06eHI0O
Oyc//nbnmxWHrmwZIpXE4YCe4vlqtXBfRavOXEADRAW9VRkowor7T3Tf9VL5nX0y9LuMYwFyVdoF
qta9IwXlaL+pNgplgTOFleleWrUvvXZKzj+zFZNAYz7hTpb3/pc7TdCtQap5JPq2nmuhnP5Acw+y
9vpk3Sonb3XEM+RqfJ9uo2wTLMSPPhNYwc88vxjjmZ68MioKfzVDI8o5zLduZ66+d07dG6Oj9XNi
7cochusXq+S7IzzaPxnuGmWp09Lej+0ksGtILAzNK1d7dZWcaWApHRN2rmVebNfjErGmba4Au6dD
E+uQsYuJmEWv4QPE51aV8RI7S6QIq1t+785TQPd5oknjwFhXlA6d0wYwjjQs0X+jdURpt4vIr9mf
qyocBcwAEb115f6J6yTpUvcfjbxq5sPp8HatoxkoMl3z6KnQEdcNNtP/UzyoLLQMGV2yhyfAxiNf
B1N2S0PknTQN9hfmtbm9KQ+p6HhT5OYFZLzK1LP8wautQpr9H6aIyUaEVZIBfsHTXMPEn5Z9G8Tk
NCxeZZuNtjt22aIdlGx1rvDdu9yR2KhvhbzIAwJoQajYHYWV0o1aHZiu37m9Mxn1JBnHtQlt8TO9
cBXKlp1+hSSgnxLTaz/7D1yvQ8g2Zw9D9Q+siMc7vy3MkdaPnyk+UWR3QYdJtZpbzxNtYtoIB1Um
zsJSvzvUKuZH7Fp3YxKGoSQcf5y+OuO2bGeJ9elMQAA12gaCetlyx3NJpBYjygheLoDrBbiPUGpB
9kzO6YvyRZSW1VEAdJBpNw8fA12Ql3KCjTdcu1hcrR1xJeJTkDdhykWXijYDU9cZnvBe2TnTL8rs
BAOW6Q1OMU7i0gNH8PB6xDQzk2vMX3YoC1prfG4pxJFRgjQakX0anB+Xlnq+FOe9PQBUSRKb5rXj
bfT3l90EsWnDQKr6cLKos9duZ2+fhVIhaWukZORPaMK3TKOMVpMwqQ1nPa7U7QtE+JGOMwmCFWww
+P/OVLcQXPPUL+8KV5nVtfxvBQef1V7NaKrOJOTRv/lZ2KmDmiPWqL9TD+688+VJTgrLPnji64In
5QnD8ojyG+BcyEl9H5F9iDukxD4GrjkpwNrWwExgMxx05/D7nxzYQYg14I9f1Rf1qG4jFQk0iw5E
AwYuF/lGdD2ut4VDCVLGiwQJi4prDSYpYkZSWxQm5H2qYTkcFlvJXy6/jLOvmzDkvIiBXxcLnIa2
UIBHqdeF5TlSJSMwkl1Mzo5zAW2dGodsTtRo9kKFIzRZ4osuHkTvRHgCPmbcWHfzViJYX0/goa2D
WOzp5MnvCZ3KmNGRFJlnxeIdUab6NcpZzlNM97+vhk+480jx7fZ6aobUzFE5JGgEmJtH8KhAdmVU
YNeNezCKQpWRLXXlXs9f6yaDyE0geA8gDtXNUC28XVR48pNy5JlpIwQxvEMKY95B6IHp+Tvv/4D5
WV+xhlpoXq0+jAGaL0qss/CcNuVhC1ISiBaiUmUjjMXsh5n5XR7+jH0pNv1oLQfSt7s5MRkilj9W
Rs2AJjnJ0XQyKBRp/ye4uAAkHjcIxNHeK3Y6Pg5tDlxrO83grIeQ8g9Bp65v/G86vlqcN6pL6Wpd
toV+8/WJSJKwUYjUdPw/IdP0QHsxfPDWMCSUeqtecsIroxwn5LVkj0gJr3WusVnT04p4HcpvEWEG
uOYXlF5oYkhhFg0c9VZ25bg+fudvV5+6oJy0FbrUE2vp7lINawiLBSmrBNZ4L1/gvKEzuKT6rLYN
xyDaYANBirvurdRrpw/80jcv4/DVvAj2+Jtu3L+TzsUZlUlaNkgd4JChDJ0e8ofOD0Q/hlnCaUGp
6po=
`protect end_protected
