-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ReAG39WWcVu4BlGc+h3tuugGeTzB5tNjTonWR3AqT1AH4+Vxl8bub/65fC045NXZ1Gb88XeIPxau
MX6XHYR/FCXPLK5/ZSUUZV5KdynZLzQH8XLTWsXduuFzfhBZ0x9d1EkIMybUqI+8E70+3mtsOxQA
Errtl/NUaunxehuPvz/eqflv12cOKvXpETMMkfVmuZX9Ixbjv7WPAO696SoPyPiA5CnVrV+v4ccy
tk3MgyL0BpgJ1gmCgPak0dklrPAlaLprrU3j1nikYvDau/SUf4u+IKGrvpP4WWba54nmll7V+Y3y
LLTVVzxrzTxSACIxM17KxeVWlU54cquQYv60PA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 44064)
`protect data_block
hwIvQtMFrSlpQ0PqMJLZbt/5CDolpOim8a2fjFBe+jOxgQowEc3FgyaNKoZprnAJpXNdlNtYAG6j
85Ovg7ph2c5de6cIL2Umy+B+XfYy/I6Es/E6Iu4L8/MOfYlt82siAyW4uVrUCGO+PTf6cIelWuM4
bRma1JBwB4BZlZHNhAOs7XQtAFBYvnovbD4Icb813mlL7gpvVykRTlHr8Kq9akPKYyyC6HJpV+XR
MO5ZcujaGZ2cYkMTLaStXkEm17uwtgHnIJiRG+O0T4F3CfSQ8A5Zbedeo5bCKFhHSABir6AWrYNR
Xd2Kp07C9zYIGOJy99NhlStD6ABDjp3VK9asg7oVStjRGMh/72Mkj7UFLxvW+O5keBk7oG1TT8X8
JuOvpuiIpI/th0AqJwuU9/Czw8N/ExqAf7PBAxIdLCwEHRE/mURzKIWCag4jl0QGt1k4clu5qgBR
p9C26RPrLwut4SvucAXjBvnmyObLWwlNd7iJ9y/ZLUjEDeDd6yugVoMvexQamtzecXbxm+T2tGtF
soFP+mNP5hTg+FdFy5HfMS6xv7u1ipkHKv+pD0xUXEE9TLf9M1xkDA48/Q7mwCObxn7++uz+HJsX
aF9mZSCUPUWER0ivfANGn1GoPujpbedEzOEbnZB7O9dbHlq3XouRI7I3uUb+fsPVBZ2fUlTh+Nsa
o0Fe8AfNDPbrxsB3jUcMutAHuMXMTbyrDl9TpS5Ywhq5sFs4FUG1/0Fbt0Jk4Bs2pOcL8kxFvfMO
6nG4Dg51O1sbpbpwwcfNH0jFGY2ArungJQc8IcdlKRdgFbwIiZuCiumlqDR95Kuv2Tf9spsWuNIw
uq5ru5WZQ36Ta4JcKwnwdC55A6Jswq18HCdMvhlxGbIU3nl+IqOIjaDC5Ei6IkmQPYbJEksb4H4O
O6ICDdLu99YU2dVHAsKMmxyZ2n/uM+G5De/wEEnbCpri/AIZae2tFok8ZWwED5XVit8HVu033tte
ZNN6kxsaBskYMnxKn9AaqZEgH0yklStRd2MhCafD+j2y8XSGHz+TpKiMG2mlh/OMpcMBP3RcFaqv
nOF1zXRsNl/n2zsWBIjp2kRjc8xo/aUfKZbPLKgTJKARQGHnTgnlUXl27IhhJ3gv6Tv9Fi7t97op
+prlt22PMv8eV0La7hoO7SKeV/IBsIHd8eTiRW5oxfIua8+ODamfat48LFatTMYqCU4sIOlBFxIW
RsUybbmZGYfu2gNP68uc9jTSdRsjipODMzi6FFvB0dGXDr70ezuf/LQDMXT0PlOZExWJs+yo9wd6
KORLWonlOmj/RjIP725Jf3v5jY0Kxjf2Or4FeLThSkuuW5lRqAi4bhjWgqJm2gKxYeb3VbyBQnUy
IeiSOmGQzElCq25BEMaCGs4e2dorvvPndm7pDnkql3YEpBI8sA4dSfvq0N1xmLw2B71/EvC/9ybr
h6ooORnHiNSkX2aheL8862PrNLdXnlWQpGYSF2+a2oyRbsLZwk3XcrSNanAC7aaz0PVHhf6vBMJd
pHITZYu0FyREswK1fcGHhvP0lA/1QMN9ieYoz78wm/7iRmGyo9PUzpprEgc5rPqlHI4mva5Y6K3J
9Ua8f7mB7vVsAs78i9XtVKJloqEncd7Z68EonhqzDkvJxoX1AguYDBzfuEawNqYhY0s3bJhfjIze
64C9+zXTGJlrT6rUOjoR7gg3LHSHlbLGpqfG55s0JHKAPhM0egkG8sH/bzCP5MT2z+cQsW6rPuh3
sofX2twAzi4eigw7vgFC2XKUxpfBC0b+nOzhMYHzNlK/E4oalG7fR5LsHr1z+B7L3dIM9S+SDUpN
JfLn+uewINZDZtW9C7yTPpvA2AURKTIiTm66hJV4mBWP2n+aCiBo6xT2XR1+cE+hbSY9yuEzvQ14
S8h/HFsrYt+arVdhnC3woNc76o67CPuNvGdCcK5ChMa6RgoAbO/NLu38gj05yudrXGT5k3hiiGBJ
+QDxzMyA6hqo1kMsCiZcBmNkhVHcWM4fyNCXV/osP3PVPnP3Dkc47wVb6m/a3FQ++wtRRYgPiWKw
q9CXydU5Sju+7zKJWY4vpJTj3JIMjOGau3oFYrzGsu4NI/P+Fu/WjVccsP4c8jvzdPa2MrhbR6Wi
uJPNHAwNOQaqFM5ahzp62IcSX0UuJvil2XYx50wib5mS9sPg/PZ4OJDYSCKHjtHRb3Ohd49Op/Zg
9ijAOJiTP3ZK24o8xVhdJFkEREm0tkuEAtEpioKDtiIS5u4STvc4DlkQIReXAmtsnnZ+rOSZj+0c
pA6rHcBx/8mKlIxLk1zywz0b3prLQ0UEe4B4Z6cf5E3Q6F0o7QSIE/BVlvrnV66DYy/omG1AEb6I
db2ptvnHu91xOKVDToYfk/A/IS/r9CZ2NAunsrwrGNRtfhPCxm1V3qQhlXBKPAu+AvQU1aGLG3JL
DI5xUwXOnms+577US2mwdiJIPAUu3+e3qD/vsJaLj5LqpwgkM+sXFdgurBLEzPGtMUagD9l1DuEB
Noij6ZU2SEP/jJLDYH6xu6KPCiFEXwOy/zfMveV1mc6qwtZQOmwnhgwGKKbvsHoN543W63YbpEo9
oWLVScK50HSTAzadlJ3x4Kzxn2giMAxG6jwEL3v5gbA90wVx47SgfMPp0+blxDyQjkKCLyMrOjvv
rSUAJJeGfAJiMq/qaUalLPD1LtRj7LkJSm/lcMOMFaUBr78FI29vKhPXmk/MtJkm5BV178Rf8P4b
2RYmiG1tJEiHgVqewbTXRDrC1tHtplpsueasQt9/Jl6CvXRwn7qZzhJw7z7p6i3riof6Xhfwvt0e
cr3UcHPLcwguYMVHgVsfRIGiLEd14Alt0jVJJ/1ElUz3OCaIuu07/S/knt4koA7FcnkYTbGz/t8s
GYee1LWt3Vn9L8RzMtIHE789BOVlu6rMW2fxMoOYXBfJADd+Wt5uiszofFB/FsQO601TQXuRG6vY
zp32yOgKhkAA5bVm+OzpYy9kPL9RleIU5iOL4Quirc7YGfTeSdjh6VMhO6lkE+eHf0NHVaHN1Skg
fIA4BqBjba1YXoanU0FwK+W73DSs/6/ZAToTgfvEFk8b6ae2ctU3l6JOroZn69tIYzyZOipO5mgq
C2P3RjrSil5+2nEwaIS4pk8twX52HL+cFgvR/5vSClWcR+AI3uh12qlLqSm6/ou9Yj/d2cF4Pcmo
faXBVzhP/Q/Xou/vM2knKA9pWo2CYyfhCgOy2crCSK5lvG0SZQA+gh1D/kEr5muQPWiN7Uh5H48/
8gSSdNnWvF/+CVgQmUNJhxq8EusMC6lIRremEYJMJffbV77II0VuWrQIiaNt33l1Bqmxbvz2Fg9C
owVldY9LF0cry1hSZ4cdu0saAjdURE2nrWUC6QRRUEyoWdxE85XvrOFi++IVd9EKCIIFoOjeDGL0
8gdPyAvkrVZyP92zpiwfBhzYe57YneOHCCrIiT7Q+DsEesukI/gjJ7pxb4NVeN163CGwfsPEFNUy
69hbgW3lPw+RbRA4qwWEIf1JxGjVcZVKFhkxPZ6UUuuYSLrP66FdUcGSLbkiS1E7aqspbO02lIYV
Y+xW14e2JcODnUn1ehvA9zMIGlp41F2ediyZkIu25GuA1LwWG0AwuL5bHDZNwdSrsrH9VgoDGWk+
xyUbmT0bwKgvcCHF38xuQDSaBlXAu4OkWxtfPwPtmy+2vMlOzUIFQ/NkG4qJeX3NYUh0hIk2kGKX
cgnc+H1Zd0N4LP1VI/rM2clhWExkUydb0GitYb6AS1bbdizQm+MMfgfbh5sGjIl3aS2zgbro4BiY
3+8RquZCroqe/5uF8P35qEcLRkksxqIB2gcAYtHDwiDXmrnPwbzmIQI5O/9ozNsQq8Xl9QePABCq
lYjBW/ZqfR8Gv2fNbzxHLsOxjE/HyHn7bSDFpBYq7D6iOxVQD3INYGBBgW78BlMq0EpAWlTSIJy/
tnT/6oGVFabs7kX9WsVYqdNC3xIxvGP26M3TWNFhLYKc3E4L9KZyM9y6xZR1/drJwSE5jsVmfxeW
TiKHoGhf5BONT4L9uGCog9VqKzuUCXUpPCq5eX6BBJRAOaG+MtTEKaETmWHMHs1zeJq5P3YhuYx3
fhVnjirvnFJkPSRvBBisQy/jeFmssSERY6VAeWrcvmjRvwZAWwfOm9NYrtn/OPk6Qo7qIvqAWLfr
NoJkv9X0ojpZ/z5LRTJhLvH+OAo6t/r3rwoiLuM+73tP6MAxA06rPIdVHx40pNht7IqVUHNdQ3sY
5aqUTqcZ4ArNXgie4OmcRPXJCurtivaFPe9wkZsv1b/RhV9nKNLnGTU3HOXQmIbw7lxpQ4XDfF6z
MGg/XBQ+67rmAedARrWBPaCzizaJ+x2v3IhhOsEjHsD0ZmdSxTxUYoF6kDGIx2an5dUExm0/GE1V
TF7Fuj4LvgtL2ZhzYR0BQRgCXCUG1Y86QpBWvSlbSi11Z2rdfTugQ8ic6LNSYSeBXTiJdiIMTZcB
leJKNjyd7ku+F0RxlqSPaFB9BfITyRGAJjMfQeZOtCmoak75267CoFgZ5OO7cRn/JVwtKRjm61Pz
6ghAWH4Aep4goGhjEhDKEk5MRAe5evvIP/nbx2FXscfL+/LHdak5u/HYGf3cAJvnSKV/0T52JQdL
+Y/Lcvw28YlnGDXNTo3ugQT/vkVD8AVH0MaPtfyTw4+BUbyBYK1RdUajLvTJRAQXIB7S8WmCuulC
EMm+CgZfpYG/Y5fzDOPH0KlDo6kpETuqxjVwOTINtS5wJvhg2iot70vQZOrPpH/+2nZkoKoNFVK0
BFNXhIgGc/S4ldHRpfoCVds6l/LN+cMfi3pgxmtipma+2/b0QeliNEbHWiZO9Y+wfzd29il6u7cy
mPGP69K2JX1RjIQGq5vKQc+g7lSecQOxQ9/BOVC5tEekb100klOhkjxz1rmWcMaCDOVlr+MZU6lF
etVMgpuw9Gojh9fIela0C4aM0Nk2J5QsFwn4U3T031uaSJ8DKk2ISCQ+TFNnCLb8DZnWUxAXaUbQ
EZ2Dng5nDhcqnu/js9Q6dH6MJEwo3zg10cisBre0/T658Lwo2qrqtpge9+BLgn5jZJLplCHYWCE1
QzVmycFnpQ8asMv6FYuhKkZy/ZIkfGCxGbV+RwNwESlRB3fPPSb4xbF3KAPxCL4jX27AnR6KPKsW
HdGBDurY+QOWqhJTdRMOgTwQCWTUB2EqSyfto6T/ei+wpLTodsimUD1GkqrwEejLdNCrDji8yFTx
fCi2xM3VbSQpFINNZZx4e/G+TAudt3fjJg4cPU0XBU3zxsMdKPdgK4OUX7LupatYSKPlWoUUwr06
u34Gu6oWYs8ENvGn2aq7NEQYqHlxWmuxpmS0dS1AnTBr5sAlbn4TOjQWiD+2wil+L6m0mZ9inJ7m
AVOaABFE9lB5kegHpdAVrHkXG7lMlwcA0G5XKMGqme4UWXZvMUcUsuuP3sB5Rqt23rauE0KCwzTf
YI8Zn3hFR/gjG4432hjZbYqBAhQOLQLokguoD/x4M4MGVz8rihIKJkorIA+73e4IS9kvIjLFJf2w
Xq+62i3yfExarifAffUyXbjzeevRJADxoaWEghVeZFc/QLHPj9WtDnyprTM4jTx7ABuO8T6Ucswm
5FpfGOYAlMCXUYUQWyZiyctccgI28zqU0L9ttL9bfZCme6HzfxxNSNYFAnQBIFxkDVhiNucEU8yu
ckMYi+vsesXi3b7L1ybT8gPEtq0rL7dmMQzeFG1Kt1Cg4vSG/Ib8oQx+l10BE8KgQE9UNAauIbGd
qVnYG21HTqdE6hpEqXJJ3/qkoaeNBFUzMCRaX4Wk0GzalGoaFmYOjtTVHxGKHjlipEhj7DhrG2hg
jKtJnBJeeU/4MqnxXuqQcmMzoxyT9pG89/pMkeXJ87+RBDiZvIGIMsJURBM8cSjCPYU+6iwNMkRE
p0fbpmhHSAW618kRWZhuI0FlIzEN+kFlv3SKJ3VMCv1FsJVXwBVohpjhpUXQAPy3cbO2cjowhn6g
1hOyrETk161MAfZIKJxEd74MTxXl+zFzt9m9W5/UYSDGuYDF9lfOsdWycN1I5BjRaDx3I0f1jVEs
cLrYv5WBrGgoHFARmqsDXN4x1jCT4p9bWdRSUMhw80onfkq315T/GNpfCLOHkzWGhfpb4vom4Nnh
dc70hz8kXlzfBQj8MG+3nX+Ogs8sTB9ikVK/1HE1rT2c33Wzocu0MT+6408EZ/Dp985NFGxg992r
z0bMq3TiCJ2dScZqRKb+4ZCil6XqGL3Sy+Gtomk5BzcZSFS6g6PSq1flG5SSf/YZqnLwYg0GzRER
bGJwSyC8x/eVmfwdo4RS+LIGnsuIv/VTqFNddH3siP9rQD0U4W4Gk6gQbmlok65dEsrwsrqCm4io
sUnJ0+gDqgAkfXbnYC/s/yXUvgt2Kr0OoYkVwSNeuoVwEuvQ4YgqwRv7PspD2t9g7985Urk6C81b
rhjSDmcTj7UR0GeCzSSK0DPW5G0mqdMyNANF0up7HFaG0dPyY6ZpOBSXfSBDZUQVaZYMhlRgILcX
MiEyVmGP/VSI4ZIvSxwVdKU9nf3paP8KLwrLapZYBwHikTQ6jK9LYOvgI9CzutmTvQMBGCxkMgfB
BLhArtE448rMd73dyqTk2uimAXdlL0j4YFutMwmbkSPMdFdElgViiBWupXma2CLPLvfOWao+dhjF
p74NeVPOzQaXu77R2mDyLab58aGgwja9Yqmosv59uYB2LobGhIJS1M/mL37sjF0Z9qcQR+2SrPn2
MitP5bCwswFd03e+VSKmZJjcHXBeUZKdJxn/47ho5ZJYSuxxHYNhfWM0mHmpUpeDQkSJH1BX9xT/
HaaSFYJEVlOjELppC3nddOiqHdd6iKNFapmvzesQryzxAKKk020DLIbaXFWigQTKjo44XGyxT8ts
7QrVqvRObx9M5NC2lwTrAa03T6VRW1T3RM4I3ZDgvlS0rqRnYzhMhhEhE/8nmx7ICOtuJoFkGs0n
LvmO5GFYIcL/UinMY8XBSivGrgI23QguNnV+yneyi8aYHNz6iZ1rA6n6zeXnCGI3pAOl8xrm/t68
MSSwpB5L7meeZq94moob1SI5zgS9t/FAmkFB85SiBkkEJ68AHOKhj9CMxrTgn4SHZJknSvrPp/uv
pvQuB6W93yZITndPKqUtjYAwfBkioSbb5d8IoBv7U2/j+cAe1hkv2K/V9RbDzBMrfUhtVHK02tMU
STsD+dBLevcTXp8qrRS0XHltXhktJ3GhfhFvSRMyZih8afV5yEHOvAIqbsDz5P3NG8i7UAubUL9i
gKG2oCes4T6cMnLn+Kcqcuesaqp97USjNTIw25IHRXHd6eyXtPDp+t/E1pbAFxfhLmCR4pTMUsTV
WtSqoY0q8abdosh3sypR/kxxcCcWIqeyCSpmVtuCkUms6WVxC+ABOPQEBXdChYge5STDeQC4FoVE
o6s7A8LntN1kG/ULm3uQO2GVBunrLLWNbgxg8MyH+AcKSfMcBQAMvEEMAcTJ16SI80WwN7ZkjhJl
mBM3Y6alC8gBPUQkElAszG7ilOQMU8y+pBEqPqu+85n8+u8YH3ShHK055JlNyS/e7p5Hmve/96q8
S02gkmZHeryh0rCJpampIodGAsMAo/20ap8L4ZPumfom6tSZnue2aJ+/IPAON5S7qDPAcKq2vGcB
mLuw1Sw4a8MCqLlRSh418pRKKUbfmP1781KmqZrKEaC/ZJoLkQRVMDHoODXjgnAylbPeIv+obNPM
c2SGdrCAgaweQcjLELJEMxBzHGretE5e6QUC8JlIFejmbEUtvi6fWemQAt9GVom71n4/ED+Gv0u8
E+llutyTy+GHsjCSZQ8C3+Os4GhM0y/cZiTcht0g7qZ/Yfi15zONFGFbxnU5kTDYLx+cmye73rdW
UFrqmr+tdKOqQCxkUyNvuAfcoP9I1FCsHgV+S8ZcSy8eyjkN1PLgrtVu7dolVbJWgbZbrPClk+Np
H+toxkh9U3UFflaU/9JC5I/vUCn6G/cXEwoOcCoYRd1L/vcYxK0gZSkmicC+F4BmMGR9kqrKfheM
XQFqJ4s1nb0QPYlADjuMCLwNwHV/3/Gf5vWf4sna89uHTm6QXBVvlyaLSMr27Nj6RzMgCbJj11Tc
b4f/FFBZ4Y63nLzGY/smnmtUlmt0868HwXvJ0rbCJJ0QhwHiMU3l0vyS9Gn8azXmcTkPEqPKt6Yq
TuRS5uUDzniR28t5EToz/1jaV3Y/vY/tSWccTNEJTUWqWY4dtjduHhwhmXhU2+ckxKrqy6Ci8e1g
EIxML9Wh6zjoKIRhekBLuK8WIOUH5KiQUfLmzSBwoT5Ihv5n5xiXxrJBdS5Lmo3rbuQOhw1cj9TB
Y3jjP4PIwToUUIgCeH87hnDip/xEKQECSW+qlkOIq3pWBNXpeFWpAl3FrBRgzbPw4liXy4lUYAPg
Uosk3CkfnK0TlyL8Jxm7g8d2AWGuGUr1XXfvGACyMbOasdQvqWdUhafurBc9ptR3851NmklY/f+p
5YICHYGQITt8prdlYk+m7SDbnlvyl8q9amkysdCGKvrSJQgJ4gxL+iLJa8U31cCaYfNnLchAAzgW
RIatUcF4tLD3/7LBODhBU5SppXg/SPDCgn88RJHqR3INoizgS5BjypF+QndErA9Xp+ifYIHgkUHa
IQ+W1QlIe4i5e4X9oefdhzhH9zk5IgGLangezzgliLdg/97axtQuAdpbhGOUU/8BSzQv0wRJafsZ
GtOBOSYW3slUA1RUoSTJ8X3JvmRwg1vHPYKycqIlmT7dG8q+osp/lSDEtMh9JQEm3BTJznn1W2rY
+OCDdlJJVQOtlUGX1QZP6wMmoZcmjeuPEhlD1J3lOFMrVhQEN4ix+uqs822KJBkf8jIYv//zY7xo
KXU6DPTWR707de+SQMKDeULDmggYp4W53NZw2VZ1S47AfZmAv8gQ3gNVKTQFEXUDL3e4/ZN8JFgF
s6GN5RoiTjk7KnbvIderFCAp3zQrIWlibgByQ297BFhV4Sxv9usFkFRAmj2+SVFTpBUV5f4yFF2V
9p1bYCmhO9grcPnjIbjfspEJbYcM2QTQiNYI8vaqegJwRiD2D2VV5y9NyuWMe5NAMpUTe8RQ230A
Fdu4rIc8T+Yqhs5CXg2IGcjPjGDy2k5BAEMd0Pk3/lSGokA6hxEAG2MCHCFU83ovyTW0ub8RZ6Mw
o3aGb2tSKH1hFvZ5slJyNX89bVUIUKQ02yfN09qXZZC6U8We4jfZ2bRnp6c377Y1sJnGcGpXo+NA
7omd7gff9q61XWdnHTeYg5cqTzPVoxNJpszaaTaBKYY7a9Jbrwx4t3MWUt3jM7MJX95xq6WwQ6wM
vL9zLXhfvAxK2cZ5IMmCm05C7pYvDERmH5Y2uNIEqHMTv992okvvHaEkzw6gWkxFwZyj9qL3QM5Q
WwS25RgCMTMegYLDoaRP51Tbk/9bjN7f03Vn9ObEyhF2R4Ny7IZcuhADqYfYy8kIRerTYf04IcNI
8Psl6HlJ0Y9P0jyjGOf8lNs07tP7l9nHiwEYNh6nJMVq+jyDe3wWExQlS8/WWkY4PwptQFYMXvfl
kfIpwiZBpDll/+yOaiDUqnXeqMYs5Sw9/6GBzCp+LVW6B2bWRH//2gA6NOkliYfRb+F7muopTgcK
RCWDqDM5wEn7IOCn4Yt1aHLVl9WMnPU2b5tZQkNgGAuHdKIdWkrhiwAeVqJbv9va+n00caoU/+gC
6zPn0ph/D5bm9C4T9piU4JWTPRtEBxIi0ikBtNU+nwundRGScIwCrNJh1x6BxiTZa4a1ZfJ0GtAq
anQwdm9Z9CPxPGh2BU1oMxyySGN6x0VoryFJa6GLut3DHXW4sBZ2j24c02HyUJthAOTpS5aWFEya
tCl14n8meSaxBHDj0o6ORBRCTqkfWzIgE207lTI+uUn8RIeGtAmuagyo5QOsCna0znfbJ8uMFI8T
wP/UCU1RUk3smpxMthnuur5m/mFBmFnH2UtUrn7czntWvQQ04n+xb4YL235T9ZziKEsg2dIT8+7J
Bb9jznM/zIdudLnP9oSUTNgf4zByo4GHFQ4p/2WQ9Zf9gXVe/TWVAW4TX/uuJugcnWZoE7QEGOSi
ZL84DwG8rj0aOTnR1L4ROEAAFEzLee6b0uqvBaN80RULDUDGUUQIbFGnf2HIgCrCrtEvvnx8lD6b
lXtvoaXO9MvCvTNj5ykdvtONHTgw1DGDIWvZ3Yt0VIX02sIrAZRkyg6FdKS9wPsg+5oyT1ZYThOT
qUypA/TkXANzsVb22cBYSRJe1kmHepyXEhGvRoxJf4oXpIajKwrN5PL2hGj2sY1NBpmh45cR44DY
pYnI9gTvFDegbSMgTWEF7ueBpD2mQpZy7VtumJnVNL7+NRi+D7dcFmF0nYSECbJeWr+pveEBRb7X
UvqiPxlTfd9FynRcBKG/CUFvlal3L7OOEzHdS7Q3EcFJw5PJYRmZdG5FZMgw2/CFF1dANrU03VSL
Xbdf1Pwo23tBYjDb80hCdivv/HhDMnrYjsboN/l/HGFZ7VFzZbmytcbU3/U2/ft7sIEjA6CwS2lZ
6k1YNHmwYfWJOvyGHJMIKKbu1RM4eFeAC3PxhdDqI+oUzIcUgFbcQvAaMO0MfFAzR3ZkPMy4Ivkq
MTqP04F44a6+wLptYnYrVB/IPW0jvF4ri/Kqbkwnpep1pBwBMcWGOOosIR4UGtSgEC4k0s/4pbgE
qhjYhlUiBlL5YlIdhwsa/JO/HXMlBZTB4qWw4wA6POHH8McoWqAU/DpadKrATkhdnvsM4PoZfv9X
UPu+tClj5peVslhkr5kgPnwifWZLJKd01iBoa+R+09p2BLS1HBGv5CyOkey2eEtyETFETDK1nADe
WGMP84ywsBWSMSMsug/fVpt1CcYFNMCxYzWmydJb/IDVJunn2oksCwxo3NTQf+yvr3m0VoTqSXWA
kWGGfOsAP54XQ13nZeUUw14xYmN6UfEvTZgU9MfdznDuf8jdnmQdj/ihkXf/7K80psKPFqfc2J6u
+e8OuwE9I2MOmKaP0JBKn9RM3ZWyhV5l9hVNcAPD8HYQ0i8fQkXndqFyssYzpNPghkjlJQlAIKnD
vnCxTBY6+n4/h32LWKVn0eIqKTNv4iyYHgEP82oGRaRjwcSviudScgzxHEFbSP/9Hq+j/oad0AiX
audZNY1YGapFDiRSNO1/ueKwSB5u3/3j9scf8zCUQpDNGroWSl367Uoi+Dy+wqI+s5syVZ9tDbRI
BGnzs4ZPxeb0a1e48HbXtk/uZG3CfEhmWYqQ0ykAATc5eHrxsH1GSOMlmEaQlbXCfZo1e60Oni45
tzLLVL1AebdcDe42i/2BCNZY66HJwr2PE022DGtM9vclDbDvAhPVAyQJn7c6Nhpg9aAH/w7zrloi
Im1hP0G6hu+pjHT5p29WjjwWmnT8L1TEF46J6u7rYFnuZLaP34/0uTFGOK2cMtMVkc+2/P4vzdRZ
jgvjuYKtw/LaDVrYkrBl4n8VPqWLYRSnjtZg+oRprbZ8LUSfpwOiKHeVYfML3Q3QLX+x7AY/p2g+
qh3EK6DUJdnICF9uFcpwErkrH5ocw9gCdLIUEI26sDoIvkJDzeFb0o2vZ6kjfvQ99zcowMphqkO9
2Sw0rq1was8BqG6l50o7Oc8SQ3iBpdXDZigaBpq3Q3+qOOwq0skoTbdEQ8s7H9ShBRRejRMC0rC0
URZzr0y96ZSAYqOn3llFo00mutXpEqCQ1EiJOmSls2s9cvTdyEa5WCu/GpSYjVijRPQu6kq4jN55
IiQRGX304wniRAsoBN/rEUI9sPBRjVIQucQcFo3NAdyejN0URakZdExvYq14A5SQyA9XOyZyGOxu
A8NpdfvkL4yVvW9Hlervtr730/KlpAHhJXb/kwREEyQajh6kdCQV1xQHTlv9vqJE+HU9CCassPW5
kq3IbUUuwVxd6qbJYKOl+7YkVXVU3qNjzr0SBclUm4akr2yYlrepvuc5B457JFYvzS1RFS8220ZJ
cSJ8YYLZe6YRBirVD3sDUS9TDb8A8Ugr7FF1VnxkphB+NO6Hiq/rimi5W/fHHT9I/4k8Z58TnsY2
RqDC2/JalgudbgZlsMwen3vyU96hiFiIbk61O91KvRJxgfuv5IJJnZXhejSC0HyX2/AcSTmwuyUS
efPh2LNUXspiV/X0P5sf3GASgdG+qBO31jBHiU3p4FeKWYisC+YEu/q4UM0go+aZnnrVnShofnA4
fbNVJqwims9zeYr5oeltYvirY0EbC32UMT105AauSE/LX/FRlsP5w1H/Y6zInrqPhPE7ecAay/NK
nzJ0K+Y6M9WrRlAU4696h6gJlX7rsWW6R1YGdracZ0RV/tc+eAvh6QGg+rpeL8YLrJIY2/lBdBCQ
c0I0LW+hUAc73aOogYgJEoXhJMtyN+nhx4UjjR1j5HtsnaWgknx0ibL+clNasVoAL/lxpC6W7M0r
1IoDDXoeo8MMXwllqk8laTlCHDP6x2esIPn5hgztmft1ZpAZbM4JxwRNQdlsvQJUrWnT7nK2b8ZC
WEVnxKDcUtHEEmY6nhrPkVTf3aK8iw5tsrgmphymMUrq1B/esjjbsV9oV+nK5n+ZdSit4QwcysPJ
JX57unU09fTj+K3zxGwHTckzX4IdOUyC77RatCZSpK26N9XU3iLfQrBxc4DCJlWl9NroLs5hnGsV
8Lh3MXNidctg9TQEbJjvidOgEfMcWfN2NcsueCs+a2gBRa2U2vQXyfAxlQwgB77rKJnTIOKHovkk
tUo8ED14YW4KcRmloJGiXi3iRttT38C+MVgfr2JcRnLg5W5RNwS9R35YMPFLdQHBqS7D328EjGkJ
iuhmI0Ir+C5BcGw/h3Q7EYXyLO9oqCuMXLIyy+i+V6N9mvcqXMdN4cr2/J6Q0YAHjVugKfdPfXoR
B3DECYpoYy/+hEjvTOBj6VWlT4p9Dm1W1uyPfpHLjfOtryaI98SvxUOMdIORWRUO6+0nDqQdc918
B3mmwpfTKFyTl2pfJxZDLWjfYMGlVTHYFF/IhfjwBpAcshL3+reTu9se/tdOVZ6AaJUTOqA65ArX
nZprYpfHR7FMrlK8G1OVfYccraQEUFcTiZnoI3KyroNCFSh0MD9HFFXkRoWtrTC9eDMJJivRLS37
m5albtXsXj2d9QrBzbMSoqTNVpjBM3dqTXcGExB+s5FqQueRTSnVbLN0nFIZCgqNt2dAxP8iQsNo
ZkurBsvm4951SNznbweOVJ8/ITDvYS5MglTjgpweJQmnwguV2+0xD/0FwdjqQ6U8nIzx4Rc+pORe
Cocq9CS8s9Y26XE9eRImG17z+A+7YEyG6wpn4EgFcjWWhPo7Ka7FZqWQ856xLpofupT0o1hXBpPe
PujQ8nJjhZRcC/Y3LVoHTclKJ4aizQVNTB2MEUHaMtI3AvOQt1vbOJEe2dO1hw0rgV42aggn7xSb
YaAotTTyFJqxpUjFqiCIjBCfo13ONTmcVLkzdPu/ZszlHLUl/FbkpwSdy8tEXNhFxyoN0FiIUM9U
twKt6hqd+I2SA/QIFpCjobc7pxHOfSpPbOZmy6/9TROQhLi0QLHoDaycYzmxWH3/quGyB2tA7jPn
VrsSFn6ANs5GVHM7qvfsQILrJRdroxYKDKZ/iVcf0YF4Nwv5NbxLB5VWVengFLxvz+OP24uhVZcz
APcUZHS5K04rq5+R/anlG3dX8fg+DZCH5KeIC3bmOVAyeHMJaHS0y9gVjrTd+/NsCP6qFASCSeQf
CpXnxvMJmcNsaeUuNOHreeOWsNIiIzc9QVwJtzOselGXYVyzbfYAqGxoANvS8MSDe041M6uBVmY2
+vRGut1CuHYy31DUD8XwIZqigQeDVSIc1n8lQeGJ4MD3e+nAinOOCRl/qX4iG21k33dkyoJaluMa
aNof2JYhHObhORcjz3d3jRLWTwrbajX7TdBcAkAuOZyIuav056VNZ/E9CYSbwgcefukA2SK064ed
pN3uemwzyRuE+DQqYXoqcPWgFKFhDL2txvpFOZdioGOqrmLimTJVvRqtx3v1UM0cllohFdcq+QOq
5r4kanGT7hrqkUrmAaURR4eiesFWDh8TlcMuG/Xb2GL0qIBFIC3bp5uHqzYzHXK8rhtPXY5qpbsf
xmjHi5SOaAuNSFLaxJA/XCDlEdwFBJaAvAiRptSHd2CyRgvZHnpQVHQ/iVKscrmuudguYeNx1FMs
I1LZJuGyX64lRBfvX7T+kTB8WPZFeTElcu+rmMZ+12krQF2qTKP/dVSbmXUlljjheah9KKF3Pz1s
4wdmJTW8cc//Idn1qCkGFXxqWXK3+qXJWc2haWzgzqPuVusKsGW1VaHKY6h3P6CSSggbJ9OwamxW
pQLNRTkmAApg+oiT0xfQLJVggc645v3KXTKFOj8hMhc3sS9As1UpTyNFyD8aVe0K58Z6KkS5ibt6
//+8vT9FwdqubvkpSA1yYkOZXV3yCzIWM+QM/n1gYmyrHHVRq1ATPIoa0RKbL1V8C0W94demLvRG
gzOgsZ92pBCiO3T8K94rui4TABKQNSJQo7rQ5xjhVAir/SkV4jH/tCI0aL8MR53E0z6xA81xOw17
BqWaRKNall3IRRzGJK8gzB5jtmE1At0flWkr5dIO3FhDUAv9zoM8ip6YdM1GElTN5r4TvCuDlVOX
qEAgW4Ni9Ki1c9/uJc5EgY1k5WtSOPWHK+SLO8FTcW8hXHvS4+dgKt+xwD1P8YT6Wq56Zv9IEYrV
DBdrzYvgWmH9SPcrmmzLnfbMn5SKs9xzNmPy6IKVlV9Pmwzg+AEDpZ+6D8vovP9B0Yq4S4uZMIlE
MI1AvkoVaaIvxy+ykBbe20CIOovun/rQgfQgCUKGhJrObB0uMWJmLkEQALUDdGiFe+w6ych4HqlW
qLu6qAzihKxD8mbi+liSR076i+TyDeCU5Lf4cSYVgExTi2wsXPmyAWVywRzUHC2gZO4QtQS2K17E
2J5r8MuJt+TCmwaxC58AaqrsjUjSaKx8b34I4DUYjns2BnYkCO9ldieYwPzBfSvmSgJipgvwZMN8
ciez2KJeuk7lkRmvgY7Kyd/OrI3bFG7ejskF1FAcw4PYn2Zs8E65NrhD84LidTrqQXMfHrY+9wv1
J0BN73zJ0tu9D0O7W2PW/q9hEf7accUUz3GBpj4XCO6ElSHhqDw1bRjhbhcp4cAchTwkxkWEF9vb
LTkCAyfs5ZWjcX0itMYrHn6UJEku/U/nIZpeigs/tzXslFf98ySLnq8h9zxPeYPCq60Cjcs1/Gwy
y/XnhaiySBCdKvXpxFcIviN6T85bi1rZXxEsKLzfD3SvihdzMvjHWYHGPBPkmdwgafnjTzY7HaQg
tNnDEJro3QrNqrgdmDlft7L6GzYhfeVZonEOVmhQjuOXApqS1Obgz0gMn1e+ZETORo+ifKDFv2I7
jOD6zmrP6EAjPEJEENs0HoX7xAQ+g8oNPthob84d+qzJe6U+gwATXV1pGqQ5LIdzAmUousZ4XH2H
MYY1Tlm6u2pwc6fITf90gJ3sl+dDYyHSpNzD9shQtU2XKAIQFcqMtW6zXLhQNDR9f4g3eXXKJxe1
7Bx1oHJj9fUMQqxoDhhTSppytyHKGj0xWT+QzbrscXDR/Bf4gfZmiS4fFVbXvDLh0N5QkS/wVSvF
sYTYmQeLl489w4rftgPoxkma79wfz6gaw+Jp0gZKGLaHxafxAgohIwCePRo20E2zijkSyv5co7lv
Qf1NO64Fb5LK/IY+hPYt7hlivVyeibJA/5HwHVtd5zUReqgiEssu7gSS7d6bYjl/G5RMrofPdKOf
dgM5ilq2UT8ckcNChF7zw/vuc/A68fHhRQAn2WTE3EBoeX/Xsi5Oc//Olbx9Pjdo1dwd6f9EeziC
FzuR6GPitEIfeoCctD155VnT2CkRF+yPcxR918FQrdVV1k6zS1KkFgVwHuD+H094V3PUjF6UiOV3
ZbzAv+mY3vTSt4zv7cZ461MknuDrtEBe0D69LKJM9rhkX+LNouDK9SBMp5hj62/58QE92mQVeYZm
WlyaoGtpsGpw8ZQNTjDgd0BvQEmtd12JHbCUSz4QgGNfE+RR2W1m8Q63vA2jCnbVPSqgQMuY98ED
ZPSmTQdG9rrreWFomzBrIYhQ31+EsZvc51Y3z2k/3siuatLErhfjgRO20MguUlX5WyWPh/kyPETC
ruUFV1GFphiBch6Ux5IGb1kQ9wv6qtTrgDQNAElZ91vXCXCtFp3n3fwjvRX9ghYS5qDp025c9hJL
p7cNjv87ynv0y4GJdidWVj9Dm6RJaUWBoYn1YsahxCY2oyN2/dvUCJ4b7grJfaTfz3fuK/AnB4KL
RYweH3u+Cb+w+0vVTDOsn7wHHMOxkwX0epVmtXGvFfnkKM879R7j8wwMFwfi5JgUe2vns/DZRnn2
0XqxkeB2SzRMcE5s8pb0SNjbkMryNEOkbyW3WeAzBRdWL0z+eJoSjpfr3rbAIg9DeHxgORbB0Rki
genVGRI62bWNRvBkkj3S5TWLhiYJLmSB4okdf9jgeSIQme4plEgGWdsDXkkRN1tJT++41u43Xaic
g6lruNjZenTQ0epiELmuglqA8MyLj0MA9i4I4WSjyYV7E/nqDEHx+Cwc70cRm8l5gULucJvq3JIp
cZSgbRmuzr6mIa7nR13IyZNyRLL1Q8o8kOv2xkbJ822UMNvrNW50kj12AZkYXjbvu21c7rKeCFj9
vaGjnihXsK8S8reHv7s7DrKSPIMOOdUvEsYLJsDxC5l08S4uvxnPFjr2okGw/WOHUGWwppYfNILN
N8OPnWOpyGCUuo6N/hPQOYL4x9reJYq4MarboyEE3qpsJXQWtAzECQZW4shQV2ECFvQpOAmmUiWV
FjreEz4+M71FyVPVbECkXURY8MidYqgDyXw+DZHwTBvzUYdzCob3l6PPH7ap4U+WvO+E0/y0WzAK
HiJrB//o89msUbidjE4oVTPjESPTn/nl2zKj7v66hA4RNsAft6eyqAk3XHYLgm48WX+kXxJFJUyn
oz+7mtDSsA/rzMSNJGcwGAIw5VkB+sBk0x0E+etxaUnB6vfdGvcD1RESMNyn8PmqSm1vrJQVvRqQ
m+JAZpy/Wdw29WLHzI6TeJZrMy2Fx8BC8gbGqBPPB5/5rbcrp4QRgcYiHyGKBDdEuZNcFUT+0+SW
c+HWqRRLHzRiNbr8+R9vHAh9PFshIqB6pS7exqc1ysEuF8pT5SBDCJ5bqaHxK26bz3OuwkR4453V
jP3Oz+eJLFaSqGmpV0cQ7208C5zh6i66GlxMa49jhnNe73y3PxnhZFfquTuHJNnvDKZFEvJkqem+
iWUQ4Xc8oSWDfBwNBtXzEYqfUu2t3jE/sfyf4p0Caffcz7vnehu3g+m6uiW0/iijlfEVVlCHAItt
WTpciQR2byB+moS5q17bJAwfOEktR2087yaB0DSa7ECkb5rFjCbJsOS/46t93RMUUi/6SV10xvDB
cOtuxiWJwNPpCU4d+ha2gV/Nkh8LbNfnDxWfqEXUyPXQixDgkj6qIDQjcG9wxDalVpRyyBSnU/+5
qPn+k98ylJQ9PnFoJUtJlaurn7EDSydQLPvf57dgOIMQdgCepmZDtRgqNBT1yCvS/HbdG1liVDW5
i/NAxpQX0XHCTtk2wqx/GmHNw/0WCLnEOrcgAbRuVk5lVK9CxiVYU5H/Gc9+zgJhuRzNISNikY3o
wcW3/MnYVhkGJugc8tQl83ym4hni+0zKD7EDObPqs6Z9CKevqnRZq+cjv+80RRzLchrbXTLq1aCV
tVllI3/hI0MQHWadRihPE/0T3hhhz8TaHPT7x49kw0YIkbzRa1tBqoxr6E1g6Rs6rQtlGU7SdSjh
C8wvS7rlzCguhkIcqi8Z1V+qne2mG3K2+0Esb6Gzqth8GkWz4Ma1om5lr+/kuWkhXONjhB7knJxL
OIFEvxrGApGKwjBPSONCOBzdvhijqpEDd1RFtVgd+5ALi9wZbHzVlGpVPbNxajnDyJdG83GzeBNH
mjHSZzfAcUe4aoi9JTxrh+WWuUffk2tKUDIiJnuZ7RSkb5PmSSop59I/Eib1rDjDrM6lqSwJeNIv
ln8ydtsdpszK85MEhH1LZFxRmG1dJiOaY7QV/aXy8kMXtP7MghadBMJKfyiJa9EdjrQZe1+kIhxP
jUMEUxt2KFP+pFBDK1BEuKMU8Rg34uCdHdgCJgzSnUS8aq8RhyBAqlluWtgqA4UJu8J8bfrHeh4d
td+PuNeaGzbEYDAvYhmTbE6tXJZrDWkij/939tmQomZIojVv7Y8gx4jVNZ7EOEOfM29PzvamRVCU
ZKC6K+uvMskwPQa0V0NRdgy4K+GT6kQ2tyN/DjVrGW6WsjwA2rKN4ihNhJ7cMVdhyWVts7XrYOoy
LgrlZBTZ98xPTqWYLUBdCMlU0vdGUgp9NorU/YHeVDtXpe+QVDz8XsEtpQn+4tg0bSvuKcpIQYkb
40ZlnUTg9BzLPHZjb1npayeFrum8EaFJjBaDJ4LZN8IOg0WQRTdJpGDmI4ICdd55YU57fM9ujObD
dwm6jiHCMpx6rAiTxAadMwurDu2knFYgWSWeXi9wIP1kRVtX8KUoS4q89xtEdY/nDpBr09MGhPra
Em3gK8WfQp+OAV9uosQTIX+CWYk+38DU0Fr+Ohk7VfMqlXoX9fCSMqTEW77IIGwW5laz+5520q2T
qxFnhAewMUB88kkcvwUfF+wtNP2uxj4pdh9Djd88M9FTM86pD1UpZDw2LkM2Naq1YDdP/pPtEuBo
VL7HIN0JACrGE11HntgyYlvkHLuJoY8clwnXmIUI1biDCp4UWSwkn+Tfr0AmznmoRjqKje64BQFy
ZW3BJTVBdHrmpAQbuAXGnCwdwKZ6y1DWhooG1d7DidnZRCJ83kmClqEFYKL3DXRV5Wzth2nDkvr4
S1E/4PoLnKUFtExfKRSWG6RiUHV+THnM4evO5g9t/R8tu59C9XfoA7xRSIUW05BQL3INZi49nSwu
OgnneuY0mA/pkeO2q1oelYN6NCpU19YVmjOWDlszFzgeRrCvw0+AfiEg6UyazGRDNF12ATRER5bN
jX3waSMPsLsD/k0GLIJCWlSJ1G0Wn4UzRTukN0frewWuUKg6ZQH890PM2FbJKh6rjA9rhv+nuoEL
G1FrOfBadO0dC7v2uIv4ubksQ2Mv0O0nYmi7J57a+JazYXp+5s5RyZURVeGE7KoAKcXm2Q3yHDca
VhzZUDkg3G+T/7seaKF6Mp/tGSqlb7rMnZNArVz3Su/UExgPjnsZBvFe72at5RtCwymqQQpx2lHi
U4gkABGhppydn4IZFtMBzNiwT877rS1tZrJfSs72cqbuQXS9KWoibMTutLXCq6NdUIbcnbIdZtMg
dJrvy1WiSDbGEFLxi2Um3Yqdj+L+Nly+sKRZM0jytsI9kpnvNcOQ9JH4usp3REZE3QTcJRlKuXPj
ekuC7YMVDtWhSaDvk1+oqimgFnJN4OeU0d7dXoo8o8tg0aq1BFzqXQAYOrtetmcRwVpYvKprYvsD
e7AMmMKfQm68CYYMsFTb68A0Ai8ujA1X8u3SVO4WTQa+nB5ELa/CmjXvEgyMRIuEVJLzmzhxjfvg
BYalqaLMIm9tID6D+VCDmT4YGD/PNET34MBm0Atkns5DW77Go4xkMyW/NPeoankptKPFlNtb1DPV
tkubEugRjeMwOvLp0L1e8JvB8u0SjdbllHM9hXqO+Hqgss8cUdWaTiqdjhokm5K9oCTYH9r/SwCq
vagANgs03qa6gOU/JeAz3/QMseB7dwsw1b/KkD0D3q/y5hpS4n3qftDYdkYXS3O+Fr+DfW5bJT82
1polt0ffntObAwvw4pEsM9tJ1IiQ0mTGKspAw6HlC1B0uB28f0iUtGaqej5cMVJcIuQ/SKDJbV/l
M1/uqqVcnZIJt01kHUg8cO7S5rqxQwd4vYhmRIhX2scbItbPIo04Pub6eGbtCXiClpeLVKZQ+VZH
UaoRZmnv9bs8/gof4h191lq8BYrtQsiLYUd+HI7tVUGHDbVLO6jp/UwONH7OIlsi65daC75f3zZ6
N/tCeBCD5EkDEAuOCnEz0FSjRvBjo9wyCR3bUQES2uQEAAlWCLdqcmHDBWm2XSLAs1OzLtFCkLmy
2MFgl6umBnuQ2n2QcQh0tRyLtU2fyzDi40Hl9d8hsq02Edcit3lbypsSVIBhgCcv3rOxcuMJ+qgF
jpHxn7kOBoPvMU9OZUyKwacXfU5cFjySs2Ff6ag1Sl8k4myh5tubLg5RY5SHPhXuNc26MnG8XA23
ib4oXaOSrvrVcjJYuzBD3+cqmIYgDF7SHSOEZSm95XfskV00c8DAfqzDYy/dC9Hzk1XqYOfcrDcW
+UeQnKCSUEEuD2A0kAzyykQZwKgHQFF5QMYZiNhZsOuyu6Kvp6/TAnPUecazIdYcf9dZWco67aCT
/9EbXtMVytwcXMtB6RsYycZmWKu3VA7qc6ja1rlr2g1n/4Io9YY1EhSoOCtxdb6mEa/Rs7EmZcrO
zo/HeHh5G6aa5o2poo7K1e43u+x7Nj+vWk/r31i0GmjdtQ9tfH5+kccALuyzsMUqSDqfM2Bc6r4g
FLQRvBCe5WbCAVGK5YxnQ1cnnSxNMQhHLfBxbZnoo+ltwKaLRV4E8TkoWPqlSkltlYHHbZ3sXPKC
Q/adfYrvcVVAHymvC1/wAELcViVxGssa1cEN7e7/dHSdB0bITgL7ct/DG7CkT7DSEHCwoLdD/+Rq
l4Ds04QcAxBrozE/02jnb4anqtzzfAALEiR7aOcoM1y7IC3REuj3jNHv/HccelslRhQsylAbIkT4
XwnU9mEeJMIw8450x9NSUBbaivWYxc694yJbGynowFpxzbR3gqgW+ojij3C2fKvMNYYv16mVcKl9
B9SHn9IUhjOZNQ4CVpxFzlmo/nu7SYh/QAsYMokEWjIBtOTGCmMWMj589J7+qXOsXUHwBYJ3vsXg
UlS7lToYyUUVN57nIpPgIE0S5LkzUo06OIKvX7ogCjlWsjXmenouDoG71cIPwlR7WEnZGh31rO2/
K6dVn1iOIfqBzhXzOD10/KKGCMFLlmlBHiBGmDXoIOEnQJ0W1xuDM7TIgYnT7EGpGt+uKxSZigrz
/0dAYmGmF3n6e7NMV3RY6w1JbygY+D5TIkWXLfflghuU/aJ7EL5xi96C5vHIvjqfLBQzV5jX5ikT
y9Jt8j4dNVHdfPNopQbYm2E6nHBeoK8LZKbFKR+za/Ppz1UreugLqWNpjouL56cIza7nfYVVHoss
4zFv3c8lwWEbMXL87qft23SMIxX5sdrPfIfuHRSTQM9Nvg2n9/4aNj+dIntzkwXBPdAL0TT7+eTf
mv1Y/coVOtN2Sr4m3aaqAU/C+t+wAqrEtqsYqTyM2W1Gg6XefM5UObBqAF+hRvRpnjats/VOZoc9
gCE5Bp8Vg8v3X45h1yhKpW24YdrG326xA3wvjpiO77oV0S6nsp4pK+Cp0kLrNziXNm26QnmcBX5e
5MpdwnBe845fkytnudJBBBQMuuGhS7utSvsd1u9h/YsZB9XD7G6GIBU6AWnsChomydLNnsE5r/j5
IMHisE4QyT/9EnpMjOwUORYY+UrXP1+B3p5GaNw25FIMU8x7eewBNNNC6u1ky6VuS8gPvFfb1yeL
2FwueZQAZwM1c3uXIXObgw3hU+k5EJqWCUQJVQksYQBMRQSHIQbH/4cYF8gSkiSuXeIxxgFYkztl
NQU4y5S3fSkgC5ci2d0Xyy/jmNXGMgpj7Ow+Jda9KaG8wHyQTr3ekFARsK6dcGJ1H0+5V3J73mQN
aGYXv3pz2oWFULiztJjW4ZeLobeuB7RsJp5EYEKDTllwR1jLOPn64pVn1Xy/yOEWP0dGDBziKfGc
7OKU3NtmWxmpJp6hYpEpHlFOQ+3OS31mdt+lpPHgF4N7BZ8WBbSLknWJQtDL39PfDuT50omYVl2l
916HEnzoPAmecFWEPeglXayVcK1x+l+Nipc2uADEqhHuKuBnlO1WUVEe+lwz8B6MG/nuOI8o+qif
GnjkI0Fr542HFM225/MHmo5UGKjIWDKjeGDaQEdAXfgQU2kd3XVe4xLA2AQiJtyMCrx84rNaYGVS
mlx7TWmfIrEAHQ6ZygUHNJ/3csCysPpOAa43Tx2MJALGry83ogOYFKf2DItVZztQdBOaGBUzs2xP
Xa29qwddJaIy+rF1ue1/1E6Y5gTlmjbwEVlKlC4GKVfavjf7DcmMwg9zY7p99dmpthqejPwNMFTn
wTu34G4dcDSYkdGlylyU3TzfMGD80mGDXgyQ4BiP1Vat7e8IdP6w0fkSTjJfm2FCuZt1JWKBt8ps
qjDTHMBnZEUG0oBbp0Ktckrpuwm5v66gI6SY8VzIiZ2hw66jRgLkLgDNcGKnNsdZaRo9iB433Ibi
LQHqVnBlC53AI1Xp/Q2ytnESBX9lYJ+gw668ForEn6ripOAdnEPQr4Xr374h2bodgbW9oy1hMMAD
c6NaKXw6iIXfYKm9zWfNdkHWcmR90iUfdqbdKXxlh7xBLnLqEpvZGQGzpsRKQq6pinnOgr9Gsxw0
lrgGhVixE53itrXg2lpQQ8lJps5cefWfK/9zqNSsQcSGmHzx0joYckr9y5D2/DMS3XFhu+mcbZRH
p3biET535Fyz7ZtpP7V83NFD40Bmr0oUmjp0wtv8XvjEHPIhn2oPSYCRaoRJ3BXqqSbF8+krmaoi
bhUHm+eVfqPwN1tLUdjevepULKqXiSJOSu6si2tQvuPxSvk/q2O5H22/aONPhcfUtEFB/Rn8oS5D
2gRSCbx3biRr6+jTc1pO+xAnXeJN7a6FMgAXGC0OvttGkqqptitlXUyzCh3dye/A7jUqYxxMTe/z
ll9TB0TeooYVyDPBB+2UVoLvYzTCCEaJUVxQyoomdi4vum997EfoE0yCmkPSh3uWe4qiZZ3+aBnI
XkiUGT9AJIPGEQOKPxbYXg6DzMlVAlAe3QM/bjfAs6Qrc4pinl9a/6nPmpcC7DRopXAingMSIk93
P9P3r8GvrofI9iOI/I1IemBRyLX+3gdvpy3D5bZd4EIciNjiLtKdyOtVXPXT+9RbCtr2Viivt9CF
lQ9hsPk/HAJoe2zTeiwt3GBCXMbI5iB1wxYF5yXV7IzNs86BIBoK9cNn4yNUt7JpVfC0YFCiVFqe
6Nuqod94RoifjbXZWWs4ppYqsZGHxaRmCtHcyC+MoHl0dOlgSh1cB47hO7jTQza8CLFehqioJ/u+
fYEprHMB9dBm9nQkPbQFabU9lTAzI2AkcyprU7gZEa9zXjfdrpnpWkqM3vwTOvAdZ8cS4kPaeYyP
5rk8ZNFZ1LFrxAPAQXVpGfNr6UHTUHR2pWF0a10tB6smgp+4Hywk9tMA+9SyoBCj8EmAmQE8sHWN
WXsvHBUvWm5no8msV0J149ut53gFm/4S3+WTkJPac3lGzHTNI0yuUp7DHHxPitiobfoyDhaAZl0D
HP2umb+udnP8TtQ2K8l0Wyl94RUWPDa7p44sEAjis0G6Lk7fY3NedYRAuLkL3zSHg9KoMN9G4qcX
ybqQAWBToCfwNg+jClqSvTef741F3+CK6Uw6cuAmiPPkBDc6jyVLN7ElCyboeMt+xfqZXp2GI63k
M3k2DuVdG4h6J3sPjm2711ZYw3n2bFmmNPKOJP76OJsN3T/qzGqyLZrI7HLu6sG5S/PBWgBYGAic
P5kEhB9QB8GnSY4kv6AjRdNlcnlq1POj3VbosI5NX+FK4BBNRFVV/isGnd3BNPKDj9bN4XEoXb7G
dPHRGRoFPhG+wKY+RgYblCU3TSqgFn8/weMi+SgdDm9r+dfDAGSXBMeyXXUqQIV/bNYajdlW0TOY
K4SRj85Ri0z4eoUdjE0dYVatdD8Y6IfZpvj9rbHFL0mQNuRT7+Gcx1KkZaQYPioBpOJtUKcAwwqr
URWwUWSZ2ztN1d6J0bAotkNrZ/WBQokYVoG9UQAtgrjR0QCf1DdEQtq6/swvFbmANmxZJ2u43rVw
Z8Be/mV354C0+S5W0WK6JXodkiTyVDyRbR0Hpnfd4Hyx5T/M+uA2vRZHUKpmQXqbeTd+nF0bzTUI
3jLZzMt5oxRJIeQNKn+vnT/TCwi2lvePTeyr0LtNEwYUxYkGbBTLvbRx83XCoS7nLoGT+/f23MrR
piWJOFLIpN58aSiP5akNc0NiEZnODydwuLOOhg4HN22w36QME/TugDTPKJDTO2xaxrtrJCt16fA0
AoKD9+qbKwbz+t4HhsaqusPlOeGcJkcgVQYWB8mbyfUXncopaOuFZqz1yrzOKiWhtp+3ucyfGCgJ
8ZvLxhm8XGdGUTYdDdXwyD80hWFa4dpOHoweFAjfPwV5DGzP4eFHGQOonNSXTFy+gweuTzovy+iX
bg1VZY1iSNEoAX5KsV+yJwH+6/6si7GmXJlgxJTYlc13x/mWuI6SNsPWtgZ2zK1TfoCYw6oYIJRl
oK/t+uBFVTSjfxHvM3AGdZ1TOGTDc4RuYho9DWuJUabAMhUZASZhbfEgxj3zkz6SV1bdW7lX6wlh
w+YKQAZKWEF/bVMN4CFEETUOZudxZGwTUy2VF/iNXE+/ES3M/tD9gaCKOSxRAegnzHQUIJLhO1M/
Uu0bmOd2GaF7uqXqNxO5Kpq95Ge0lwxXwP6yolMOmZxGLPLu2U2ZZjf7SZN3hXXqs8NpYmZXtEiH
O9eEpyI/xNpYOy33oD0z1hnNpoTsgxKY5auz86+w6tEHfxMmWdvAX0dx5CjWv5ljwBIKssONYngj
eVbcCbjGANcgepVqvRpF3C5e7YBfmK8qXvgnBjpYQFCZUzpoVAf+b6gvy9wa4qJwYXXEa3aBirUd
MPWFcY6YLjlRrscsjZXIaDMp9jyyzAmer2WuA0kBY0ea3PuYyPJ2Q0FP4maz1jxr1HFc9s9R6lPj
/PVd6CoRgpkWRdsID5vHe1pCg8eF/shhA63tmsgugIsaB9QzegxjAHBp2gILVFdgwafFPOk5xSrS
s+zW1KxHTOfqZCultQhmXP/5wHO7AhlSJAEqmIpyHHg2Emsu3hgqahCgnzod2ScxIaJuXROfJs5f
EUlQqPyl0BL6xufjFAO4L9OJ4j6Hw5hEfsqtzICHMFhkNu9q5P8bJ5erL9dDbq9pW/EIIUMn6kWw
gcUO6WPFP1nnHbN1t1hwX0J0GWbdslLCCnJS4KT/x/EmmA5IpmQ7l9D2z3MipWM134Y4aw1ujWuX
ITsneFLY+vq73t62NTpvBy0FgqHwtj0Iwn9T84bZ81h4/AUwyftQFyj+FDR6JHIOJfWPkWwju/P2
tiTrc6KAHXJCkAGucF68bGoXQ0XjmOCkRHQLJT/1f2pGprtM/n7zj75zoh+qxBPGl1gh+uSWYVQQ
S66sGG+FDBjbVXKSOjOGSKR09Y9bc0pJqO2S2n9IFW9r/nf/1QzRyRfXVhXpS3qxFAMgMQg71Uzm
2fJZljpjGT5coxULYs31WTV9JYVXbmLdVNPPpV/1pIooLYE6mP7z6pBbXJJVlSExw+u3fJ1QdEMC
A/eV2Mql20ItNxgUj3QWbr73e1YT3ueyepC/2QatKPEn/y8KE2j+xDUB0+N4vsLOhWibGadN/unx
yozJYvJmmVnzX8IA5yVJPxWnoO+WI1JAkvM/STk1lUEm2BaWKyrMPJO/B8holEc8lssHHHw7EQIL
2nJv5yBnADsyN8pPS8Lbsi+x6H7RHsJpjdMvlUDfLdawlqhfTC0vDD6lVIW3ynjfqBQT/SOG9Bc3
ErmtPTznmi8fPwvm1hyrvAiECxctWJYUvkiMAam+jsb9Z7v/ZYrL+wa3UXpwzI/4EdO/kbIjvhE1
cj6aZtzglszBR2oHBoxfqUM9qRf6zsE/DKW6y7QcZzgfe4ohHO6yPjD/EI+Twhz6ZMg2A8ynTaM3
kW0lYycvmdm0HjUJgaFDRaNqhDyr07fxlnM3q1uA7LYYI9wrUYXDRxZApNSlfBjBP8UhuuUiEJsT
cPcJzCBtVuiZajmxhTWj1gAOgISMNRrrWgsKUGVprvz/r4KsSpizFf9lakPSGyH4h4slhFz8WiRZ
/ihqANGWCQTjpb6UjG+q676f+z2cNMBqPtZAssQvjX3NYNvqZf3lBp1GvKX7Rkt61YicVFSfd9n/
BCHiq8enDc2JShZM8PXS4RGBysBHZsIcIfXoztDssNKXkim4CSJHT9oQIlS3crJl8BUuLRcCJ7V8
0hYS7nKLaqqj+jWbx18ji3ZUNbMiR/rNPYztx6Be4b61fEWu3V8FE3QDQNKaq8H9uVAd6VaShccU
bdMHIaR1wp4gVQkf/Rxl5g25vRXMferTA0wOlgSl4focgTmtluLW/kjrj1ZUIAoL4vRJzB2L3eaY
pFfljB+W/rngOND6+Kze8qy0IvlMhE07VIuAriR9rJAgCIxoggqthHQIU+T9PHr9/gKHcQTz1tk+
UnwW32oXB6y3xisCDWkJeylWkPX/fV4AiDuchg7GTBRfJMbVcEdA3yfLKqb2i5U8r56lSPH9GLl1
qKgs7ntiHIIFKoeazR4z8Wz0+x1EkDXzMgeDZ1Y+ZpJWQMci6h6QbgjXoEMOXsoGls5+e9goZvaA
PyDzwVWHXfvfQhdYTum2e1JO8WxD+nDpddxDujCK6AAQWJYWzPelT3b6oCURQAmqx2Qy1bQPZF7d
Eq+mPoWTqVrKsp6Y0sHyGhjn+TCoN0d38DXZc5yfsLUy9inWL2+aYBoSqupenAJKm1i5brGojJ1O
jhRwqakG6cZLpiFnoD4nNRP6LvDkMgtcb35NjvOgGsVEOZoRUWKlKGVUP0cgT8QVppsxyrbxUdM9
USdZHPkOE6F+lCiGKLqG75GXUmUNFn1jjarjgJwoffCamM9CrkJoLEFmZ1gcBMWOeR6/9mbwdx9x
QWUPvlPJB7KnH4P8Aws/L/p3Io1ut/u01vxU0ACjJUNKxfJ8s5wKOxJd6NZApf9I1M50iGwKbBw+
qDO0k8E4ZTPSxNgUdJ6TleOP2I/Pg+h8TV6h7H8+p8FTKoQ4H5UxXOaju3FzZSi+rgtUzjKqNq0H
vH862u00H4KjfFm7tZUabHCRTSg1GqXYbYaWZS96LVFjeix+z+MBVheyUj/pZ9vWGC9JBhm6hpno
h1z0GHEYtnHbQ80Su8AgoS71nmsK/a0kkhTOMkF8G95Hv4iRaJ/pQkeqp3Pumxh9Y6XQLZldV1TC
94gWka2CNjpRB+KZX8JyPjp5tplsVh4yd5XMWmY4RsUx9EiyB2oFBLsfsoHwWk6/f8vcwSEZa0rR
weX2YsZt/WTzQ3BzVZw8PrYtelUexNYHBA+UZ3SyOehfb4ikykQAvigueh/FGdE+bZ0znRUEum8y
Au4mskGNg3yrijbsc2++aVITf62gEZ7wVM02JrjKei1tNCw6DLcdaD2ThVKDq5HOLtfBZn0FIGa5
fzZkqnxWXLI+94jvzWepxaCm7mTFxgyrgRYl1dR4okImZUxY1/GynwsDQTcQOfU66k2dzVPF3kvv
1C/wtj0yW/IM5hzSMoerjQqIOYcAFkNcrl9nDEq3jWqPU2smeKkNkIyuEkaz8y0jDYd/8cC0p+Zo
CQYwCfMNnBC7ri2M2i+bXZkK1pg0MlCbHor9AK9ppjj0Ey4K5GQap0qPquMjyv8o3pX37JpKAZsO
0uFXUib1iYSvGY1rDu+qPdcvR8lv8LYT320TB0j1Fb1X4FxEuI9sF50cvZmjNLQdU7mqHZo9+n1a
tQ6pP3EUeXSsIOkblTgIip+C8a8ScAZvw4f2cwWtmOl0B/BxOU4XYtOK2SjPtwKpQsCBENp3uN2+
xZp2L4Q8WASQQqASyLwV327JiHgkxdI7V+mscWhEuX873HSkJP+cyNpB3sMRSLwrKImBLz2Fe09x
g54l5GPbaIk1TirtWqtXEV7wOxnOcgBJDwo4Sdf5+07f3i6fZcPPe4GHsOK/a4QNeHN+GBuMjgtS
j4DwLWjgYwPsxf/NDJK4DWmorhmFnIr3ejqGK9IhwHdSplLRYaXcTYbAr+1lQy0FiPUkqFeTuM8k
LoPNCxgvGwYuf5Y6y3Lt0sse9WlngeEdoyZeBzCo/4oe1hdoFFPsouHZxLawdfGWONuacTognBK+
evnupISwm7m2VHNKly3dJJ07jqu7G7RyoZVrk6ETjkn/wFqAnxD07QkUXjrxzaK30pigCfqzVPvq
Ec+fuwIRp9KZm4XXw+E7kwF5HmCbCBf+Eo3iXXPu8tYAnrA0SslmKinZVGJHLC+ewPw8et9r0Zze
8RL6i9BMp5e35Wjn/YQl+pgYczoFoT0+mW+OvcYTfEz8ddBt0SZfOee9PsV0gKs/nITu+5EZFYh/
5At5M0viXIe8QoMm1wO4dT58Ncyjsa0hdooq8at+RfzKTZB0USkV7z/MvZS1IFNvZ7dJqq9+kEKT
BgH4PsLTixujg8KvjnmSZ58ndXICSzqWKQfbNlO02uHSmMxtH94NLACVPt24xfA7kVyC0pSg3Wcb
I3J1JGIWApF8UGGkMZn9FVtHE+CeEr5q56m31EoJ+TvqFvNdlFJ6Y7mOE4aakTZbmtYaoAFmGf9d
f1qOa+HoQ4yxKjvsUIYV6um36Xa1xgXvtad80w1olGSiiq7QdXaq1hDSKSqnexI7EmLSLpbHQyvb
S5uk9yiGC8sUdShGa840+oKJSn6XSm4rueMKm2R1TJ6hNF4XcI8TOqnB6chCofUpUiJdu83jiQVL
uMJjaIxeCGD5owmbUT+eIWPCmL6Cy2WndFW88+QRMiBCIQwOVjSHNRApde3+hHyqj+SN2GCWTk9y
FzhlejQGe1jsgm8fFVLYStM5snmDZbH1N/cnpLi6dgdK3urXEHR6AExHW8NZYK/3+rxRNKL7/wQI
8A371hYOKsuatDgrgyDhDblQiEDKbWDeL2WIk29RU44U8qHwDA56jwD6aifIb+Lq91/yJbwvV321
mMuCEJOEoejS86wl6S8kRfVKcwphfoqYZ98WEdSVlv4EKPGuBBPYSdHSoY6ISvn8TqVtcG2Ar5iq
UcaysjRz08NoHAXaKhfvUxIOsDerXMVW56hqx/YIT0L68112vdgTBAXiq39Yu5UlUCgePjMa0U57
73dSf/H7jjJTbw6jKwv5Sk2qrVfwn0PPNaL0kxJgGAdhhXAkQQi4fo/mIJnqiT6OPOiWkYL/XV4T
miLNUHOwLoxYszAeYeK2jiYp7K8IVacmHjPccjmIZyamXqAERNXTgoXqoXXMi6B5jRLcNiiOb5jz
4rQVyIF5FrIqLuO3OTHDU5dovC5aDI1gIj+6kFfHvb0hAPZw92JsL7DMwjKvTfY/IO824dVJzQdX
asu8HTyKfgwVd7YACOZ6IsDP2Bd8NxXM4osTmpZxaolQklukM96FCVIZuIv+B4wZYlRjHpl0L9T+
DbcaCqAL4A+m/p3Mh1tn7zVjeWuqWD69UwlLgiWctqG/JfGnl4IsyNJfKiuaZxPfEk7RAstMhkuq
EWdU7tkml2uoOqlFnDNvPQmEJfQ6iG/mARtsBOMyDupCRhZ0YCYYBOCo8MhPjpfd7P64p9mj3FMa
xWRgXD1WfyeK1jclNW0zdq66StFwOF087zqtcfr559H0VTy7+ncVZO0RRGo36eU4LFxD/aXrKKcL
qWGxWwMJ6Z5MVHPpQZyYHhYh+YczY6Zv58AQojej7yot/q7CTlnjL7M+JXA2k4+/q8zuEl7HhEIl
g1Zrqc2YupxKhKaZ2WJBfETtQj0TEZ6AJ8U1EZyotLzHWHPFaHI0ZziOx97HgbaWbaEnU3Uvpr6T
ycl6wmJevlLYt8TodEokTROkdg6rftLKiqbvXyLQOXMkxz7zhS6BWTh2t8PMvz/NTxVzIKcWqnEL
Rv6TYiFobNRalUYefVQIwLpiSd5jcTJ/tF8oCryOdi3qwR6jdU2p1A18irzfxPho5eXi7WS95An+
NLi4mWifdMs3Eli9Kwz3o+DQXCFYZ4sdKlKNnfGeVk3Go7rjM7T5aZaJyoO0+i3uICRLIUWCFxC5
kH8uDE12e/5GJEF8GQqSo9dtN+eZDX7Tn0p0l8QhJglMUwlZyx4zVP611ugVOJ0tJE8UWcNcuV3q
mvmDolbd7Q6RBD7DzOxMK0Dusy4UXmQsS7VbHvYuS1KFbosqB9Ask1Cxg+o0QQ2nFbKFJAgsOxkg
SJ7XvfRRm9b/QAKnPntA8WNIKHGh2roNqsrcXe0o1K9l9yRP7nU3bD5huGIUuvbEMpNEDhuUZSr8
ACflalDR2lNCktzg6QXl6E8fuDUhi7ptO5l7QNcf/dRfWyyiu32gP83QaiQFs3smMIVyIcfk0wbT
l8ba0D1NKqKrpAOGTz6FEJMCOPE2D8iZfFOJVIwtAaDak5UvaP94N23+24lcTqfNPh0BlHDBVGrx
SyXvt700B5KxU/xr5tXY8Ffw1aG4mp5TTesgfkk/kntI4MDObEcjLZQYl/UaAOsxJ3Gb+/qjc+nD
0a13657lMfHTo79EYc9OL0FCLn7mGy7EI25mAiQRl4z4YP1D4w/wl6CIKKnIclF1CIsuaLno+/kZ
GICweAG9HDxDqMZk+bF8l0eir/o9P5Ug0PNwEifkhaQe/lgC37oacYAViApn3YL/8BmIRUNgeCpO
aTKu6+SkJ/CAybauy+EFkjOj4e2e0Tc3oPE4b6xTUYPtiDN2ulnGYIFH6AvK0spgISCtgHk1Jcig
IyiR2uBT7IESXpZ4u+XIgwjPIzh1TvIJAYgkOvENoF4bfJtxq4keOX6AGmj0IUmoA4c8pA68kVIo
wXHqCoSk9CF5gmErAEtc9Cca2w8Z6tJHoHAPfB9Io3KkMlUnu7vW6v/c2pkOM7dednqQRjKm5p20
U1Elz/y68yqvl/aWXg096p0NLtBnwo8p+tFwRkduM5+eJSaMgrVTXrm7mq+UG45WkOJ+2M4moocV
8Fa7W14jFtIKLh7Uv8+Bh7LhG0PCUCgXeFEVPOmHkX8NuKq5zBWBnVbdNyVyOf+o93tXccpXtNnR
kmBkzmuqotPaTJ67JoO6i7sKsQep1rNUR8IsZ0iVCwqzlLbPranJWfu51S2Al/7czBHCnAinot9E
L/nTiRLUrSPJxUe5iJFrdY8EAdqoR6AMX+qOe55GYYH9gRIi/OJv7hqhuFcKHbOMeXon7fnT2J3Z
lXpowsqGXLuoKDgPrQJRlNU0A6B3u2IhB9QdO8xDDUk9FvK4QA7JKY6A1W4ZEpAYge4ZHjpOuIkc
tPlM5MvUz5r5QRLr/92VyV3CU1WLDVPViJPuqGQZ8fUvHSoL3sRkAxX4HoiKc3nXScABKHiKic48
R9YY9lGdE+UHBmtW84C3tisvVv89o1gCCHhCbatA8GXcmVwuFm1mn1bpX89A13ae7S8MF//SsBZw
Otx/g2SxYtyPDwBCzy3pg6+maSVcHF4qYSAWplcQvvfLwLVNLw8Xq/k+KOE1OmAe8DXXmM4BAQa9
YEDDhvYp54I7Df/JtHiR/MpSzIE5G5a0CooAX3m/tegMN4VU/3J/lJ5Mod8kM920qvbaL447ea/U
XRLHde7JN+2iVebHJAaqiVDpUSILnfZpvmlJL2dPwncakAKebekYfxKoMooN25Urw2rha7SV/seb
He3UbcgnrXsFBJQN5rLlnBSmqdjO5OO2ekTLs3jN8s62hhp2apiFKu8NmgzQPVtcr9ivZX9VXyhC
lrevrLE7vtROBXot6vHeQmTzsbliGXv9zirS6v/vGYcahBG1gLj0xuBtPPLsq0uElixA+6zNFhgW
jec9A6bw640CHqGNW+Cv1xbAHVnLJ2hp+fKsSfTfjdk1DSwf0y9yxdY4yspjBe7IRqfEd/X37+Tx
UOaSL/h+6xAOfq8EwSWVcZCNkKKI0G3Zu9F5kCqVJKlYve0MiFCi/It2FOjMR/bQsKzxCtNoGkPi
3w3smTSglZfukfvqUTxmSDk5qFRSPzypHc7c5eJtQQplsSt2ZLWEnf0kHUsRK2OgrxRzXSaeW1mO
g4tBaUdKL0l2fq23yxMOSn/Up3akpfO/DMo82Y+ARiN/7q6JMIgF1JoggYK/ACB7YTO9uTyiCbtR
/nq8CGbNlwApiduurUFu0mX4Vl+fgWE3mFd9YPn/YNn6SGJKNSg7Uqq9fEekjRg3lQSnPs2fQWyx
v9+/XxM9Q+prUixcUrLVIgZqoYBpsvmzhJjViPwkRrVE+JV38cYCZEv7GfwBPqFIbOra+kDUkdQx
g2wUqCGbntsZZ0N9YlddhhjO5RunsYtmzXSW4iCqVbGWY72qzJ1w9uNdox+Ea1eDGml+arjngPlR
ce3MBC7n5qLRBk/+7JNUz+x+H5vS9MGEPzuxIqRrtl/Dl0h7ZmNIi0TM85iXH14t9RB2KPlhKbTe
i1biOvcGT5Wv7MwfRVsiL7P5yMY+RRiQcmHWOYGOAUrusONfQJX2mkHSJdwte+BfuVQF+hNxzNuM
Jcw74LcwWHnsUjkDJ/gM7PLsz97QsYDnA+dXFqW+n4XkUtEt1NHRCV5jT3/a+ZLWPhlUPvZ3x/r7
hZVGkHC3K1T0wpYGSZ+trkhfhuRxm0FQ26YcC4Courkxr74GkAnldrpyqgBfCF1B8ZZ9VDdV4P30
FqblbzJO+LvN07rNexWqQYIlIpXd+w2d5gF83907SFDGAFAx1yti736qB8w3ZRetUHqvOPkaA8en
2PKAcn35YTXxfYKxWUIVjmYByZZug2amFCRhA+QuCOTeh8gOoz/miiNWcuwMUWRC7wz8J2mN2+PH
icw/OZRkDnsrZGDXiD77s7eOoECS/qxAiSbIny5p+FSgIFsd24SJD0dAdFEh3DOnI0wmqIWzZlkf
iGc95KrAttM633RVkC6tyM7iobfGOO3NtigAaU+NwSi1xLH3GNuuIqSyxtbZORFJ4vFE8+Msnzj9
5WTjBa609q+aeeOViJVe9MIBjT5uar5rFCpXsl+mg0FdItHhyBt6JMqCf8kWMiLKV6/f+Jh4aFC1
qOOGBVjZWJYkW+2DJkrfLekEL+ZhkFv1P+Mtiep7OogFy4tVhZsZ/JLKRoPaP0+XkTmiM5gjbQ/M
s2nOkEyXv9MFtALkIzR0zOWgXsZjgiQYB5ieGEHZdkO+/eOVycVmfhaw6np3t2kI1Ji2/y5qZOXX
YiMJZOwFqNTg3Ca8oH1tcwvNbIgpzv81dXzI54GLgEG3mqzgl/N/zENoRGWZF98DuUhk6kcJQkuz
oSZ8XbkGgO5I/e49PZTvo894nTdNlwC+9gP+c9N4nvSNLL/NjKukpucQhgVK7k8AlVIJAgCrzagn
rtZwLWroKDMFJbUyW5QNmPJzwRDBpBEWhLngc2aef4MztQMaziVWA2cz5xULHYMUlT5bpPajD7e9
72ngtiSFUpcsc5Eqjg+yWzMadrhNjFRzw8Vp1JnUXc/i9bqhl+qV3CmPK8G9ubRf8W4HGNePq5xS
HwGPGahjOHeko8AVcG32CViKE/MrRZm19NT4ZszdKaluQZzjxwl3T3oZ5Fw3G/WKBx09CH3SevtJ
b60matln5WrMXU8YIpQ9TlLjc3iMPU/9QUXhN+P+KdNQDTyvqbAG91+WDTFFeM3rG5vBVcPpUOjQ
pkD/TL0xkKspyUNYJW83ZlWAIVVXnLEzmtOzLDF+8LhEy5iTiTuzqVB9Eot1dIdZRX24zPJS0R+4
lXHwGUuIDwL85xv4S3LptpdfXmPJnilL0oGGgLKu6emH5ifLCaMDkSjx6QiHW/pOK5FYEOJ1zD9M
rctrCzaTvs/YZkmeYT/kRdhiTJFoM3Fpqk/HCATosET+QmbQGOlmfxsqcyJOTq/atS3VddF2p/mA
Sotbg77ocmsF8HAQMuU8Ct+60zLjKkg1vOI0426kLo6pdVkw9mOUCdx6LojNEo8xr/eRV5qKOCuA
ViAzr7X08gkliIwY0xJvLHaXAspBxi/8eAVA6+1UteMgOSepS3M20sCB3JFSDeep9vAdsjg+N98g
tibKWBuTPuxXfZtSOtAU8gi+Oen/zv+IiTXIckpYVBpDYlIgHgVJpvTDQS2Whn1gzEAZquNfIOVV
E/a5B/mF7A4fDSE/E3IsYw1wnG6Jr4/84gVKwLdYPDt0e+EGfSNEsDXNkE8K5iGCX9M9BU2emaNf
gWLso/zvdrhWbDe4IZjaiuYH6oBzxAh5dbMHJSVEZl02oGoxdtulagYM/R7XNLhpVmNQ8gUZo3c9
7PDsE5KVuDyq7MoZY+sxfrYAke/DGIpwtZ+O4AwpDiR+acxp1vfynTKHzHMBbBHI8R+HE+k3beQW
eRzvz7ce0g/ssG7uDffVL51g/+9yAK84crwBGkkimP5sS99YSyG9jT0rfup9ZZ9fEuSA6Ggb/LFH
fetUNAWNc9PymBSPZpaiupNj4rOU050DkhAulRovysokXu8s9MRQFwon4yjqmMsened04fPpSPaP
9Bukxq21aZMo/qzXtwfmEaTqhAMMnF7PbF9LyIQ+wtRRFrES8lsYz13uCKJ7hBOIil+cO1mxI+gX
+evzwVgfOrWjG7ahEfNhkEyZMVhGUb9ZNrzyk/TCbKEOOprM+ZWJkxtWQMwwoRQ3AU21h+GLdNMJ
LDfmxMzd2mIJrLKW3PetkJkqGqw+uu0YM6pwm+OrjPCASxvxQKpmxTCJ74ji5/hI8vX5PBdd2jJ2
ExhOAMJpFmQ9hu1BsEW0OeaPz6ys04ASjrX3ubikvzCN4vb5Vm2bh1SVjBpen3E8pFdtU6f3ETcD
7dAudSpEJfeYDfkxbZKv4Kib+hOwX60F4MdsrSPl3tZpzYFEK4+Z8je0IFYEoRgzeo5PWUgUNAz1
l+jA47rYnvCxJCRIQt9m3SB43W74J5nxN2y2WxZQZI+StoDQBlMTnDvix5h65l8e2cp7bf0MwdCI
rM8UqAGM7CSVaYaShOKoNDJXW56diYUDtItYdhhoqkHt4GSn01JWYopgNMtJY7x1vNv4CT8m96Sx
J2GTl+Zayjw4VS5M2Qq0W6p4HkKxs8pbjfiVKH5CHb+xHs0S+5G1eHjrZRq1QrZ/aSYzGynkm8F+
LOStUYMNQnJuxSXUo5PrD41J9BqgZcxxYazSaP6kXGab60S+tuILpxhYSQq0oTpNuQPrHfgKv5R6
ovDsiY1SySHA50GrhxL1L+V/U1GRfeMnh2GCDoncj2pmA6vDISOBxlKY3NTJhudLdJK/8oOvjdci
KPn1oQs8xcHGg787ww62VRC2R33gAlR4wSdDnPDCYY5c/JxKQupBkgpijQKvBvVABEk18wvbzrQ5
yOc+vZKQc4bCBV5eVsgd2vOdR+RB7cqK4ZO03LsENWz6+lyxYBKxffdpwDp1CiWE0r5oIp+t8LS3
ajQAx19Ch33adkaCwwWu4v9Tm/uFg0lorvKHvogtgdTqJi8OZbWLCLgk/nvLkICJlDhqgn0Cu8UU
cWnmwEq4SbXjq+tXkmwYxA3R2snrj2XzLZ1Wf72SL5UPrGCMkPLDJMA38mNiBNejGxrk4AWmtzFl
Mhbt+gC+RcldymKEtLuWcL94ToNsAazQ80+ZXSRvj3b087twX4uPZLepIa4dco/GeDUIEdnxXFHA
BZcNzMRj46nOjXcNrZ6jz0rLhNFr2wAXFPkCPbPDjj207V176bxiMlbDedxLhgaZspgQEdpx5chA
RZH063jwZ+7jfR7r58NSrBoJXhE4XBBlfbXDdRalp7HqG+Wiq8+BcKmSwEdTIJYv/VqPDRZ43gKM
eHiqyOHTfnOGrkEBdDYacvusHBmSTd01rvUX9Ui+0Bm0c4QX05UjN0jmhPrxI1UlxzKNSwLYy95v
GI/THvNs3STDQqWcNszrggaAVI43ky8Qw84iqypooCfQ5RPNzHRG9xZY1sQRBq5xRsoLeddwPmJV
57N31xSKmPOfJs4KRzEw5cML66lROBBkNXZNqcMc32HX/aXNU++x6Y4+brHosc+Dz3zzuhBttiPd
qzfFAXK0HhVxsrczYdVNyL+ukUlDW2vw5t4VkY/eQbGPTEf8jdtTDSedpmmmqcHn6uai4LLPsbHV
51H9qukklfT+J4fsYj/rQJZDMXAZfgn2oTaZ8MVpILTjS2B3gNephug1YXAFp/eHSIUPt+vLaxEt
bU8pfX2uKcfF9MNEG0ScYRS34OpXA61Tg6DoNRjBSdaZHfs7qpujlRx9xmFSIY0u3pjO0M08epru
QSCaWEN8UwW9MbdInrpP0ZMGzz/Tky5eDVlDJpF9ZiK7ZA033ztHwm/lw70ADwCaLGG8bAXysjcb
at+8WaDqp76coFmHISmNLAiWkfSthoIy2I9vV81VNgbJGObLCTPMg/4QWqb4u+uvnIOmG3e9yjkw
EMrngsMDNtFmvnOe+l/mdETNg+Z1SdSugzTYbdnHdic+lTV4EIxM/Y6BqfkwgWVex9k6dlqCXL7V
Tv06PqLACwBn9Y8lFhieWThVUuzgX6pJlBz5lsK+isnmSHCETOlAcUXZFcsxaw2Vu6wJKkuqJNLR
Sxekswyqo5ZKNHYuGa9VTAD3TwgFWcHwumaKZaC7meP7O2RDKhpvk/LOQObZBix05TikJtgVIr0b
BCNXuNHnCxT7iFZfk+Kvt2/Vd6vPXjsHatrf9sji6TF9ul+Wi2hGjRzKvzZPOjODR4qF8qQSS/Lr
Gbvx/NSDpLJ4nWMYmE177UNVjHUtPpjOR5GCVJLgSlm6sjsqLJ8xYaMfIWMNVXRkdI706RnTX1ws
4He1rglv9sfyMFJBBAt0pknOIZ3trPHhelS8KPjWh5K/ADBWOuFOm+6Zu05Ut2HVuI5wRZ4eVc2D
0Xkx7LaKS5eEtbQtHZSe9wge3ERE1JnKdmwGzx+/NkLLoT5OSlnNMCszCs3Egsje2wp0dsdwPdoB
jBQXyWlzXXg4JEJNPwjBhrK7gkIfYv2OB4hfWUGorhm+m19xj9a46hM+Oi7LH2itQQs6uvnBK7b3
p0FBdwq11yFvycnpyVE2h2f/v9ofOaRD6ArSuZvUQziTC9mf5pnxKKg+oobk88qxEkUOeSfGAzSy
I1EX2xLtB4IfTjh+ywlxxZeen+X2o0oUJEu3ViS29h6Aj5rpJNxy6nrg0qMpJU3x7F4T7EJZ15Vg
nNxiVgWZNw0ORR7La20ctTl9WW+Z3gmu4Y+bHQSQQhxxWdFddjFFH69sFOgSI5JYmSOzbAEmbApo
ONLUP5xk9J1GritSlwhPvz8eHZMeCaaxyPcpPt07sEoPfBkmga5g6lZO6vpyA8DpO/xr/U7Niljl
Ph/LhTNzgTxIB27KN1G8EcnMnMbvZ2B56wazUjt6VgLcLWd/CTjwaWR6yTPPwiXh81rI8etSsODb
UPWDam6oqISI+DyD8RDGNasci0xEi7BKbI4zwfwdH/7WpOAX5vf5i9QUbxcn8+vg79sImXqWPr94
9GCJKJkY47fXIedruDvItd78enVkMps0pvaqHJvamUVS/Uzm6D5fuXLf5mRylSIj9zyp8loSx1zE
pxbipZJVb7szQ+H0dpr2PGh09o4ihr/DLTBUTz+HxiUxwIdcAN95bIbGG392KBGwW96ADkr4X7pl
RFnGStjoV/v5esThgOph1pa+lzsQUXU/fYJNlR10YGABoLtJrba6I2qyg/9cuVnLLE+0s5QlPMEh
NaCDo+XVhckqz1zmaz6wOecio4h7dEGRfP8QOdMza+wxFHAUUFFCF8tQS4KeQ7iVr/mD1DseVHsj
NN1l9FijO+eFfwJB+V7u8ui0uTFnMcxaxprlzQas7Q+Muj166NOaprqKl35PlD5N85ep9Lxe4g7c
no6m39MwdomWYVY0Hb2rvnnCLwa+2xLPGSA/5EOVwW8WG/rvgmCXDpRDnOqaXSz8xruA7EfotMpq
m5Bv94lXmLfU+WLmlrZtvRuEyNs8gOHiwnmATVkevm90kyNcpnpa+oC+jU7/FIDmWJb87gOmQ8y6
ZOSFmDzbygQBf7vYvt6B6wOAgtwzx+riDDi6vR4UKDFBg1stQyKuvzLOdP7wOTh5uWwEjQln5FvD
/KadZxAA5gJbW3n6X3G/YWFlhY/Z5wgSWkcHx63awX2DZOOlg+R0/v+O6t+RI7NdOK/8XDyF/IC0
rpKO/G6Mqsx8Gb3EWZ5p43Nr+/G5J3d66z5yzAXcrDwkrSwYsrmzs6FGs9FPbmSDO/YNAKFe9ZDV
oxoU2tzGKf9rLwCXDg/ripg4ZPVwTQ7ZpNDAxwzlLcYt5CWp6iiLXf4noTag/7FzWTKEBJ//j7Ri
JN8MOuGaW3c/6Z1Z/LE0OQY7cBp/OTmFooTbLuNOC79vyCJEXkEYgWpDd6gyPVfrKnnjC4IomTug
Ry4pgc1dA0+s06oe2kepd1X+8uB3or12vgYvx9olaaores/N9NRprFYGCEIG7T3g+j9ckgth5swn
96H/uedK4DK8OEUluaTfsDDTcU6medlh8P2qamf6OZdWN//v4l0tudx5/gRPVqtdfCNYr+hxXPPx
uCXGxpGYZujkcKAb1fQNcA9VjWNqAgJKc9+FR7BWBiu5WtR4IVLQIU8luVtOwzP6EJihF3wpRT/l
j4PhJviYHJxYyAOcEs/71mbiVzWSDRbblyHEKJWGhSn51TjRPONTLUO8qAwEtpE2k09p4zBPbsk3
Xf0z57dIN89baXKFNK6RYjwA7LF0aB65aaOTpKPcIqZ9Lv9MtM0+2JrcV1SCUg8dUmYmI7rdOMpS
CtPuSTbZ9I5eiwupHrbPHxmkZOde6ka1Qt9hq+JHdUpe+2UX2kIdhiiyoCLRbC48h8SEdruGjBon
8bevEiW+w6Tzln5e4DZS+2WXLOoT4XT+eCLwALcok03+Y5M7AytlA12IGgI6DQFEI1k/FtQ9dHDs
lcOaGLo84i8/4EvZR5CVPirU/wa1U+SOdmSpIOWO6ly/Ib60uufpDKI+bEJm6ZHVaNI7ZE+VA2tp
AC5ddP0vMHJrtHslBrp5KV3XhwA7GQI4X0UdiVd5yt7S/zR3n5SIGA67GHLo2Aun9wDYKpmKLP6O
ww07xGFV/L1kpz4SFzQFTsNtfM6c+6WcXg65Zre9qQucHLMc12HFeWBZ2Faw9KjG7lxfQ8rjhbVe
nfvp6ymu/B9p0Hn19ZrgXzRrwiQtyICQgCDcBxeOqRRHfMsMk4nYVyp1+nl8I1lrPrZdSBVBHs+c
tiLIu3R4rS3n/6SJf/TKzhTdLEBkBQMThHM6jo/KjpjZ9ZpfJ3JX6rzRhuXAnab63JZ5OTpYY14n
fBvPZwgBHWh+HgXPvK1u+HBXcOiu1TyQsehg9/EOe9t0yzXvpXyfNn4TYseKj4dkkmiOd2i3s9r1
VhRHPlFjngfjyNbZgL7XXyTRJP4CYGXkdtssbsKIgVuM8CgNG86wjP0ASKSLUHH6O7Rq1XhjmgzH
wnDrd9ouRMc4QDI7CxXoiq3yinkbsBt2jFf03XG/rwDCwW3CEJDIRUdm16uxKT/g9A2uujl3wTAU
VReWScl4yY08TcbxDVyXHIuzodgPQnFFB165LkCvBjrpLI1Pbn59vJTZUUYyMBFuaC3fQXeydQ/2
8aHgJ/XYLTdij3wlKWjzLM/a/Ca/0tnnfJWM+FUTSbMtbJ4HgyHtN6PcBkClPRAtQFvOpMONhLOx
OFDsiyQnXF1KzM14/urcZmoevNMsBbKhXIGN9bY7EjFkghOygNqf+9To9tXRAPSsONAeVbrlKPmR
ue2uiXdFukoXmTs2+QuMKMPug/Z9SOR+LhPauYnsvRx2b/wfZY0wbzphfuqDHoSzIqhAaUzsPAfB
wk8tya+tDzfJygpNE7O90BRIBL7Y37Tfe/EQvfqh2nBq4MazRDcjw0rFecotrNsJ9t6T/gcN87CX
mji+hyTL2BXLDpzSrB9gOWeGGyTw3geH+5vfU4GfmGcRZvUyQxJJC04XVNhuFUrhhWuQkGVqfKWr
VzVLp98alO/TRsww3o0F4ZoYmx6okSRFJCK0bg9VLkh4ftRDuS29bQ9psYgpkB9lrpTbzm2taI3+
E8zB9AjowWF5XI48FGIMNQSVac8IVBI5V/VUrAghUGDbkYw++2V0ahPcgLhJJiokgOWm/QivezRk
gxMSHHfAgbh7Rm6VPYmVbT14fzLjYGWa2lsuwt84WRVwvVVguCqrrUJ3i5Tqvr/6ETvELSWEIiDL
0R8h49CIUmlBDOTVlUEyF2i4XNV6+2sF/wkOX7xgAT2SioyV5DqDsyLBAE0Awok7Zne7Gs+tsjqd
a5ZTs+FjkIJa9DJEnDzWrtd9GD+zueSy1KAqpU7q9wGAKOGBzBCzIMkCb0VTrZzIIygTidVZbV6k
BbHQ9AcTssbhui/Aj+KxwpC0OtX5tls42kuryOgwoQGU2s5zYrSC8iT+kEWBOPGD1jZZr1T+3Raw
bD3cZ6vSpKgMV/ONg8v31S+/kOa3axGX1OIwRwY2LD7ay979VGfJsJPoW4QoHR4EEVTWg4NBvS6d
+0bQEVxIvzk3/sgb49NPxH+s8jSL5yqdmbCSdDr7QDmFojvl0ICPcHvMsNPXeQdG3EmXsKJGA7+t
SBwbyuvFUYPFd6sWMn10wvuhUr7B6icI2W5N+82v+AvFUw+sInp0TUuU9pTuzbA7tvrIu70lzSk4
rnjmDt2r5qUtsIB3IpaTzKD82tVA+BIFU08IASK/SLwtN/gVaNmZVp6CQfC8Oe9iu7IoQCBlStfk
o1cMNE9ct1EJbDXipuUDfvc04gkrwE5e6xw0LtUIUBgO5H727vOge6YPVh/A0yaMEUkMie5BKQ2W
+LfCeqPHGgfdRSGzozEfhbV7UQVLdSSYOsfCMDr/SWI7gDuxQoA6dagcHt3zD2go+hK0nd5cyf/j
f+icTNX8Bsy558Qw8S2WSZyw6sIBB+cshRCK0vJtFw8ExgQdgZDQ1Zg7fiu4eXOMYH0ZMH/n3z1y
+PKblBiC7smpQayV6LSxDePNlzIN9AJhQx/IhwbtF893Whsn9qZFPX0Y19UyPoiaCMS9nZdfVcEr
7xYV0eln/438g30yXPbOB90ImRB+ynMfhMX/DcNxt8IJjUWxOHTuQw+XhbrCJSHNCGG0aCPqkxbW
lpvmNeNVhgemlhPZCWRafYeuBKNKZcrrSFsFNurgnFHnQc8w22UeQdRJCDux/Nq1IkM705redQSW
APL/gqMZRGdNV3NVAsAapS1ZfBFx6SZubV8qHjm1ek1KGtceKkS9eeVYQ4Uf49FZAzX+CA+U15Rb
RqRh1dBt55axwtaB3otiibzj5KLSE7TzlayG2kVOywq+eNHOyvylqP+qHeSgaIpPUrw03CfyC+Q5
o0lZchBivyLviNAHC5x6J51CdbirzuyfxuaE5xPUgWhQ/d3BNhOxIUQ2V4D3uRuvudyh//hFgdNF
wFcFqSAPGTxENncXASBbMJx++yVg3YBZYN44qRd/5TgFldoMGwOlmQAdAV48I3D4xoxQqBXHWGla
FQ9BoRBKRNesN1UbLpJzjYjL1e9l4oKTu2VQNMW7Ku6SFvkuhSG0RkNtLLqLlZJ1oG8doLPR6Jxv
Oj5SdF9G3jS4bQzclWEVqBp5wxaFwgJ685ivYeQdF9pdqQlfBNPhM9EI19XwMHt/48nH97pIMs/O
I9sRarm4RrtqIYgjwyyohPgqfIGu3PrJIKoFjGWC0mYfIVuCkk/fU9olTTTgpQU5iOZousHeWs5A
Pm56cFW579QOnzxXbsqubr04ePT8QEnm04Lm4zcA75lnUV3eA+LXCMoc/jDEfG/TmBdLE/2g0Gvr
5Q2LZlIhv4HJDTIC2p3qTauTX69fxOafbfRQvdnHuTbcuVLb69DNOdhCnlIlqtuah96mNsykZxpv
ZXc9Y6M1T38d/FCHopK+QfHkvWtS9Sz678gxSMPd8z8TyzWumzFyLhOZqmZblAEM4R0pFc5EowCM
Zw3b/fm4NlnqBXX/CDRvdZEcwh+SQp7Nj3WT6jBSPC71unmdTVZ/CbnAL58yL4HZLDsUukIJg1Oe
GLPlBYYWxnzuBDIIDH5BPBkRLlZDMijEiTLIW9HRPrwY3pjHdev7tiQYvJOOagqL6Dmlv2n7Q/id
Ggksa1fxijppE/YPbXefAlGtn+LgQ+IhmNlRY4LI5YptxK63RL3BJxVreWDJzSZgU8GImystizOj
DtWJ7VIEsXrpiJfQqz0AJFwlNrsQ5YdEdJLfm8Y9T6b5oSv4Oxlnx3j6A7tSpyaLCQCg6h9awLT7
WuvI43h67tLDQCqy+qjJYCIbF/TKbBKTy1kBxryMV9FSUvKbS07V9qwXbjMQl4MYQubtndf8sTy6
WVl6JKj6bFAYcvsBdUxzruiDk89z3DKfPl/bJTcTl+pfcvC3S4Q8IhA5RHDWWRcnIzBJVBb/mr6z
9ZK1PN/RfvjpY0tZI8KTvwXWrqZioVRRPkrVPvBzvY5B1yqs40TVqJ2h2kpNz38X9qdJ0HeUX0vS
R/Ieyy5sJGxudzc+FE17l9ZbLosKBSDfIdVn1r4s+RiaJ2sBkwWGHrpekKeOXPKvGEvNKEYv69r3
sfgKqTbD4n1Q3+U/kno8txLynDTiWmAuW4BHbvchzM3Izk+pNzOm/ESNpcnA6wcEdhlARTeGc2Cm
aStrKf7+FuoZzucD8++y/lfjsW5ud+IrPXdurdkdoha2YsARVP1B9fjCnHgAhx+rCobYGUSCTwjh
QThmy7+x7Fsf5QydVy9sc43BfpOnU8wVq9JIXgSP64fzuZIhqg5mVNTfhBMavkOT46/4zPYAiYD/
bCxo1Xb5qOSR/MI/SMFie11AKgjfbYBfjm3+Rkxp87l8pJJgoeJzWIR/r4yGRJ/ikx94dEA5fE7s
HELK6PITAC1UIpVbs/WRhP+y0OyAcBIQx7GkzGcxpCdAOonxJ75W5wc3NofzvlqYXQjmOW4WHx0O
dB2/fDqaw1pRhLlxi004X3Mrtult5EPbS+2gZitNuh+kHZnVMEnzdHDO4o4Zr6l8Lk6CJUDGi/YL
vdLBC+0JvBj+W2OESJUdVEa3Oz5nUI/wS6Pp1HzPiFJ19g8utn78E2aFTk5S6E+nx3HDfcNdE4gv
d0JMP8EhO8TFLnPneHKru0OfpoD4Kw7Bbc0LbQqQJqoWNO1lY4b5hTDxqCKIMOgGJuGBdRIutx17
F4wNQHnucoKI9YNf7Y+cVRDuGjKbKJYzwqYJgrCYQh2ZUJZHqpvPCI5Tau5/cBBFNI/xTLXY3WUD
67Mv8o39a4am/RzXxmJKAzqeuZXcKu+eSz7m49NZ/N/QcpfO5qkExZjIFhRwqgpZUvILLaSOviZh
0GnJozElNhyH7roji8q081nJYJyni9pNe52cEYqOhIRUyqMNM7eKetIpR+im2y/twsExEx4+9Owi
/yXgPUaSazpC8bbC1w0u3g3GiTJsm/JrctkBocchF2+smb8w4Ys/JY44a+HvNKVfJjjPkskr3O4u
gSv7r9nR0J31dmL4y+JwfebGBPSpjnUwbAVsd9SFcAUIe+fr4L8MhAOX1LpvfuI26GYu2cjJPb9q
UcHAXP5Q2cwOs3Vq1BfKiTp8BkSN44q8/LEaKWxvYcWRexQuOKMujQTvL+RaR920MrUqBrNBECoU
J5PzbZCuzWD/du3/CubeLwrMpN6ItvVuYlzAiAXupVKxrPyRUjosoSolN99nqGgHffxnGQNiDlFw
Z4xs0Y2l2Z2pdUGq1Uno3GVOf8uwfeghitl2Y65J+WEJ4ETdgTQ5z1SLYLGDAYiys9bVLYTHz8TA
rhzqqiU05yJygC4eCLVN3P8+AdIyrA5SoWmwV/d23AK/GNGtQdqqjQhV/3JqAE8YJKdMzsYrCBoS
sQxYw8xXEgbeJB17nDt4ciDteGldp8KPKs3Sodv3XS9mj5FCcK8+hoXLEd0WMs9nSObMre2sOGay
t4KlJi0aNYB8ijkHCslXLB4l2RAYIBqWz6mEWSPD6ZUeikvXorLkEWaMf5BYeDOdICn0GjokiBZ1
DlYZ/FT8FjtyAzgDys2cp8jiSZPjbx18GjNQHkh38tIIGBrfwb5ZegR0r4VEOtlk85BLS9VgURZh
eYMWuzVHRM6BUViWOggcGVIi5DNWAsiK33tyR7LFUkBKbU4RyARtxn+nuNGMkVHYssb4wDrvZ8Vx
DHxEiQjS89Txd2GE4NVPDVC2hksfDsRvLnvHDvoA+gQjGJtM4xWVprbo/zzOnz8a8En4wIsWoj2L
TsgZhJNrCdH1CWNSxYw3C/7jHLSabGRCV5NHn7vCokljIWcdIt+nnEIlgbBa5/O1gUYhRWTfF9H4
YAN/65gBMr2pp/fWU/yQ9yq5RPAnFvzkT4/Q+qVAdEVljsjYzUZAoUbmWW9KDPvXHdFaBfKP6iS2
woEt/nm5l6euBiK+xesnFUOvidULe9e4i76lGGxw8lNk26smh2hRjH7oVm787OH3cU/ReMhhwMoI
QFMhb3+oDgvE5vT8jAXeNUPCiY0gasMobVSVEy39oxkvc4GEPM4GReaPF2vCDqTBCIYSs6p6K/c5
nrrXm0W7uk1cK0REXqqWdksnhP3/wkZ/KUCuPH5iaY99ccBV36w2xFJN92WBa7jvbGpw0eUM/vwP
YQO5jOb4FqIJeaojuOKhA4jpMHvmjfsxwRwyTrV/XsuFAe/yl4XP0eIC9NzCNh/pf4SUHTRGj8hl
Ua+CTozB5diKPgopx+KLGKK/RBz5pKbL+HQ9rqsV2djE9yzB+2p0bOr/hkmFg+aZPj1wXDo1LT/p
UUTOWLh5uBuAiEeIbFSILo8wzVo80W0sKtkBT30fGbSR0Og4fABpqFdMccoN1Hd1F8mfnKR77Pxk
jfkkJChbVw3nL7VVsWJJE/zsvLwxbwCrIUbZm7x16KLLJGbY51KY4zlUr1BAdS8aik3t+sI7Uxzr
vi2p5eusCu2nQJ7PUFivDMJQG56i42uTe+5weBcxdUsith6QjwSdaZP4OjdZBLLCBV+1SbMy9dY+
0VfI50bsSlxYuCth8V4W/aklMNh7PhJ68I4AIXJ6+3aMe7QWJ9q+SC9KI1dtYQtpDbQh2yzTlSoo
P9VEzEGByiXO4fxaSEXSZqejyogqoGsAiZZc9UZoAV3JLCT+rELgDAC2P9ZS1vubCm33f2MlqXzq
OlHipfyU6XZ83L2RBQEjFgmlmzFwHpTuyHG7okQe6xf2Cj49QITAHsNLuedeCGEHmmfAT6oM2iMe
RDkZhaDZ2WpshPB45SVOIQ3fVLwruW+X/mhRr7CM+O4/GkCrmTXnIKnjqhQC7UmPHG72ld6Bf8bs
lkxGv5OgYZgblUhBV+VT/S3CpDcWd/AlFCJHCAcGRy3bfn9glkU0Ejfp43aKIhdUbzWTnuxKORD3
iii7X/yDCmz1Wp78TovPy2yE50R7B7BEtnzn2AGohbx4yMx2nnHkmHkyJL53OCPNHWy51N+oB+4f
waU40R9f4BNRyByD6TM+LZyNjfi1YL2MFM9jX9ZZLw3Nq54CPYv7YXrcYLNfuD6LC709uwV0i34x
G4mlkPULf0Jo5uf4bLCXtK0XWnlj8MfyYY73iXKmdsiuD73jdttlz9b7Pypaom8urCE4gkYZtJUX
Zd/7F6tfnI6IAl7GjE4AF99QselRQWJk5ZKZpf68cevGLjbAiF0pp+JM8kIFrf9fDnzf5y9GgFWX
DK+TJuD8Ac5sbQZFoWPqa01LZbgNcb6kxRV838NPIldV9tSnRPyLpsA+gGoS5SPxkAoka0pqElDO
KgwGwA2vgMWxJIu17JaarOwjox/GbgcjnKu5dywkI/6eomx/OOCqPu6Bs9tfnGPKKTiaNnlA3oJK
45KvL4UoqfxioYBckRPEpmcJJGm9amp2yb8clRfpGrMk2w71mK6OIUxOsARk0YPa+MIWlzWzcsBY
FzZc3BvAc1unxQQIztbnEM4beUYIdSsYba+VuTuBfkg1X2+94TQOsL8uvv3vbOqHNaJZ04Xmcbf/
3wG/xkzKuFqV2OTxLHDOwPUr8Cb5z6nVc1jPohdz0illEQfHY4CnB8qWswESe6+tMuE5JAIRqwli
GrSD3x1Aadkw5CjwsUJE/BehvTAyZYf3rVUGVoqRksoJDNXfQWJPjUAUGiicrq289ndCYcGKTNH5
8lB4stuoQMdRlXoQZdTbQxGycEPYAilHO/kakyMKg7tb+gHVFXI+ijuQx3nbjJjD0FESjyBCu1ir
oBcCbthSeAVYD5ThgDHnYeUwCHBburUH4b/6KPXZIQdUBdqtlmR+/TzxVlBlE+T1HtKxU7/dYGlU
RXG5HGFeaAQrVbHb7dYIKz+XqnEX36RNL9maRJMPw2QsySJ9IOFfw3RDlt9kbW5hcMXyGjboRafE
5SgCnSPfmBMVk5SKCs2VoHxK/8uvojudAsmJZrMqR04wMiZ6VAhtsA0LCF0TRJh004mcC9H4f68a
SGFTN0I+Gm2HV6r4XyrPac91sxLCYHcg8wMQmOp/PJ+EVxracLBc/QnF2ACf6X+i4/lrVCTcD01N
D/AxPY8s44VVPTfRpjgJwH/mfi1crzHHL55j2PwZQH3y9hcd0oiPP63li+hTFf+NV+peM5CatTOC
jqf/Y6YL3op1R9YhrtDC1/3kUeFTP4J6lOxhhMed23BK4wvjTjq0Kb3jbsKR0RCWUDc7pmwwQnUB
uro8fEhwbVmm5dUWUsuwoB+zxOOZVJwafzZ1UkXavq0bcMNlBR1T0wb5XTrkjvBEnDlGsVttyx1i
hvX7BWFxep8XzA5J1ee6SmWkD1TPDRCXPNyt5SRoMsgBeyoHgs37QEHvj+SLloArn8j35OHPzUUZ
OsgZEyMtAcZlXLx4TZNRAJjD/hDZbV69Kw+YthUwk0IKudNSBtxOFfNJXkI6+kCEeAMeUF/1VB3y
FBTpbVd5ttXREVsrXHxCf3Pi+7W+mwntULq6RgxFwlPA0PXtCCvgtc6bleZcxG36QtdP3b5FTqPO
zJ40eCYDjjR+Fqrl3ce4ESJJlkLysPurOZvwD+F9KY8LqkiYbRpZzyUejmMLItkwkgMYAuPLHDDH
t3YmLZ8L7a8Tfx1iMVedxOYDA3UVktdN91MKiFJGWEtBzBq07TgqyS/uSt4qIsmfFvQeJyqn9T57
LxMOvih84o8l1Br5JyNbqyVL/cwF8It42275GziXB+rIpu6fX4qruLAv/PM/lba91KQavMrtBp6N
36wGNXxR6e4IYCCPSwxxnXM9TdJKGChR9NyxA0A2/yI+r6c3yHOYA51mDq7k5ADtR4JCndDB97bD
yXZsrFjEiou9+4D2D+/SQvljwkq2a5OkccJyMbVv6tnHVJwpfSLDRCG3RBQUqNDu2/823jHd3zEf
NWWFLnk4DV7cu+rCcN2lYpub9mStOTruIh2RuAbgpYBjV2MfEB6uymFGJgVNHpZlBpWNZIlAbGXx
fIeP7pRvzB9YW3RtZ60/aof91rELt1QXaIya9DH1xjUxxCIctCKdad1MkgJcs/QjIpCguOZ0/6b7
WuHcPUVyCqrSCJXptHaqoqGgLPsCfcLeAZH4Vr7pU6Ode9gNWRKk4k+2LYwORNOzBZUP6xKj7d6c
5Y3gO8vSaCDP9/V5W+jY47nczhqCy8idVYblZeaCslKpeMgQ6jVmtOSOGX78XU5i/OEgiPXZmg0E
t4a6qb+n2DyfZQ2Bt7yE15+h4ugDfuSPQ9fmMdSc1rEq0qxYLfxcl6DLEGQMMj/0l8TLS2JTZ5o7
ybF2VYuFCd0Fs1WhVFFIyP9RcJc233SEOVyYYaTvybAJJtrkg8ziVpXzuSxBhqUSxQOUZESQN8Zd
WFmvb+vG+hLBg4YOVvZFj2xMM2Gb8mvQfh1G8C3xNMm4dthJQ1tepj4PR9RkYU7cfYRSw1kwuazN
kYNl2F9aoRfpkSGnDQ4q6SegjOgO/xehtp4DDoD4l6T9lvGjLYcF7v8qJKb+KbW0weJ/QpPeaIlb
0K+p651gIy9rSI2YO9Ff8VEC+bFRL5kxcERmhvf6LUXBqnqohWCxAtc1omAXbVsnA1rH8oLEfzwn
cOhl6MdFCtHVrdBFgKAa4o6ZXv86EpbXmZ2j8AYBcQSMnf0yuIJDk+WzNnvWaN3UEvCAJU+VVQ27
+NXWS6wftH87t8Kw9j3LSa/JVSx1cSiUMz3YtCQbypcrif0THFs+ko92nyOfYQMs3l/NBD03FXHN
5xxQ56Ifx7k7QEqAZZOTu+sdNNRwrODN6r3EqmYoFmceLD6PzUjPGwWFOFjHr5ix5g95gdeBEEAB
VcmKFaHdhZ+3Wzbs7we7DS0vpvgfxZ0xvPJ+CUNavRMHagg2+AXEPwkeAmqe8efjLs17xVMnj6Qd
3FF5bmp2eEzeZRpGDh+zcsUoMmhZJlrVeRe8JaZbqJDNn475sJooT8ubPuom0RwjhFJ5k8nfqqws
fx+UQT9bWp+zh4LunVYzn/oIBn/et6Xe16MNmCmsljsUCX+pCt8qdfyZLAc4pCo3NHjtQc6Ykw20
V+JgwqBJeFBb5astooZMxpYQexILfKt/2xfBZRZ2bKWgj4kW4BXZ3SXkLKB370Sw5iq2wfT4gwmG
qwnXAZGU9Uo0YeOdWHnQG94R0xZwxc+xlAqouaI81Yet9Qfh1VRAyvj8xH1bARG0mK1noLgc4Hp+
V2ZqqyzR8Bj+Y4HluB6Uxbjh/IMQhIM0IibY+hMDyemUckornED+wYDk5Pfv8OaZavG9YqqJL7cW
+kBPYjXjpm/9LNsuUs0VCsjpKopBKRZUYX6AwjIza/erdxX6rO2aWZJDi8lz5RryVm3E26sSfG/l
ziGH38S9M0oYNa2mOdwfTVrSbkuVXEMBhqsQD/b+qBxry/XYCGivhhi+4VHUPE5dKJyLlfLxHhqj
a1wHa+pJIvPnvza5Ive/hgihWyAHb/C4Qf24EM8wXIvSSr8dG18dYyNX6EcERQO1LzdL5Y47AHHw
pO44ccMVrj+OzRwc83EjZMRVfnqA0GURsDVcgnO1EcXkMEcJrpIEY19jwV1GfxVq88oi6HIgVZ+N
nqPhyn8rhXIzzfU8Aw8t0OCAbvBaVGiVAyhd0PncM6YMvIWNJBXC5IgXxVtY9JNDSO9FFghZ5fKh
SManr5pie3tOFfWhZbrUP84Q/bfnJXM2sV25bksUsBbQ1CabDeKQ9B7ezx576bI0wYzSpWDDiOJB
CP3xSgP/XV8bVqT+0ZeLFsiwC/EH4onVkske82i516PUzgxrTug5dvhuQ3Xa/UjKFQuufurnJ0fX
IqEIuFsBGMCGCGh1gLOQiictC5aE1u94qltDLyijnpb8D7QUlI3aRfjeUu5M2EWic4lzyUT/sS99
Q++iwg6D+l7P5LHu7nOvyVeFbL6O5jkAPGMr1/IfwM056uaRhCp/2rBjmQV6/xZWjjHV4BNugLC+
ZH459nHXhdKziBhNmL8xdGQxfwkzw2v3FUYmGlAModFuT49GS1C7CL2JKaL86zc0TwCII8TpkuIM
ABjgt+w39QI2IB3qcPp4mMRQF3yZymCuzmrMrpHfocNWzPppkHdyoPcPeLA6hajDtmBpMn4wEz2N
KKc5Gi+6tR27HqrQhsaNQSXFZAPegWOIxd5x+3nceYTRRPTxOwDbgGGqiQEiG7XvUVplX5cr7dSE
FO4qwE5/kWmAekApOhSa21Y5s9ZbX0zUujWQmfLv/KIqOib9EuAW5X+nvl6OFU/fVuTzdEYD5KGe
ppLkUmcnHlI7YIsl3s+OFxu8uGetJLYyf0F734Isaoh435MNWOkyd2y1n1QMcQEsTB4NlTdVy7ua
kkr3ondh8P2IjWadg7dwvD0oRMEp1kAiGGJ6kdkNM3i2ammv3I6R2K3IQ5/gLNO7NI09DNNp3DGp
Ae41zvWZf3ywB0wu5MeZvAweEmIy8zT4c+GNKDfUgFH3tkdg+dPhwtBgIyfdUVmbdOH0TlxzpvjQ
AyLkA2g2jajCpejSREq1wZcoCyxsSOcdwf9Q3ASL/E0ibMKjwHZmyIuDT9wZQRZZPQVPpEcDqfeW
OlLwn+OXDcnDuxxp5RmtpBpj8XBGe0+xIUSitkBekYi9VYlOorABQ8RpB6GtIP1ASltaGKc7vQmr
DDuybrM46A+x4B1ufvupq6GXoPDB9rnqx9pzJkDZ1worGKnFHLJIoP5o0kRoP54xnHSSi26v5mSt
r/fub9kTV7Z0B3Ukr8su4GajtURiuNaZtd9hfTMSGBMJ8UogainMhgSiEMvbmq72EagHc3GrizE8
VY97EZLFGk9Hblm9r12GvBJMbrLgP1F3Sz4TWlugnjnihCWT+Vfj+x1kyBfwoMQwOvHrQMBPZY9I
1n54Uf49Apa/BRrFMGAj0Vyrl2bsxZ4OVQ0CGZQw7jT4o8mG+C6sVCZX1II0Ic/AyRNtKLmfPHoa
ulJqRgjxxj3hZvUmB1/Pant0dELJjY1H3Gc4kriDV+PNQh8Pa5w/jK3wS2hZObCpb8PpUOgrRj4A
bJGdgr2hLiiC6eURC7aCRItwpKIjSVavnVK0D+9puBZ0TmnQgWUOYU3fPHoQn6T3tIy6QCYGjJFj
l+UcZPF0kVV70xoZT7+GNg1X3bWlWQI/4R+wWQFhN/sJ3bEDGckJY2mwBKdojyn0GsDNq2RTTsZ1
FGgooiH8hjCme/YQ72y9wsOttQz7kCRQnIKWucPFBBRlwllGUMRuF4N+ER65vpSJxXPq53cFDY+P
8uTFFvdblbB6rKVp+/lqAah7ndb8LCUFlQQhj9aQX39DARPdV66BAqgYYHGgME8TbaoId72W3Q2A
TK0+pcCbQPwC/r13XT992FslC8JTEEuk5GfMg6AzHY+D7t6l3fQOMmXJEumD2b/5pJ7JNCrqOZ+G
TCikekKAgwGxrBYdvC8MQinDGErFqqC/KfTbhZDsOaj6lLTY9aPqwpF58NhJbevXjAsv/PgEsZ1L
YJHnX7GlPkQRZxaA4VAzxxNGjKKoAuAuBUPZItRSZe+Djd/Q50VCxXIc+bT3Uwe5hkJChAIwsM4x
TQfVesui77mf66HWJ3yFSFaxbwEBAWW5+fJXfA+ghXGUevykGn4X3yj8PoOS52r7n6zZM/B81p5i
zxF83kJahJ8jW+MAeKMy3ONNncMN0oru+HewynFgcJlBDLcQKhAy2Ncvos7Rn2hpWxXdoPT/1nvE
Hs64+43rO8qqW+IC0v400xfpHMuU9k+YlYpmcfCYcVYG4IOjInaabK42gCAJXIaAwodT05Saqk2c
CTsoKaAfxl+3VRVtrMpseUUqvE9qRLzo63Q61f3bZvf3PA1jCJgmFwJZjjpWFT1KTmm6DLxRbWZw
MGLEQRZ4y2hZBcKrbu+iP9n6K2NYPLX6Wd2sht8u09PR0288d/Po255eJvS6XWw1iW5gbWCf7Wmq
pXTAPl2b1drJIiD/Vw4LfeIdbUfBjFuwlLev5hyKrNGPLG58OSQnE5oemiX95aE21/mvXlToPeeK
Vb1npNLwbQmyRPJ8p1mleJFc+r0Itb8oB+7K+PcFJhmwFFZr33FHG0DfO4+Yif8zce2QZ/CfS6fA
buuvFsIU68uUEOoZ6liMcVJ8PgdR50cgNLoTTZ7gcsirWVYR/TzCZspQZj1Wck/X12F/2eazEp4a
X88kSK7P9Dfg92WH9VmqGwVsWPQmqK4DGZ6kOjzm+c6CnB0wn/BpC2E9pqjOsUK4R0/fPcVXlwS3
FdJGXFFOeXqJCqFnWj4hmyB3jUXQ0i9U+RIJz8VY9FjhMDeT1hyJ3FR0TCmsk7wB8UnnR3luNyXg
ptFwYptFsYHMdlykexcm4tY0ARrsd+obO68YaXvUQFwkNKBNbmn/8MEgkrOEkeHAUCPIROSZ5VjM
OfjABQnMwe+rJEamJbEo7Uh+hkt9Strlon2r95RpF8zQmt7IuRlo5A6dM8gQBQrwDsx6iIQoAFoQ
npk9mvKpfI8EU3EDykAQHfAJV2pEawYAQhEZiDPDuyblL9ivdvDo7jSKKZuyHvjSqA77BQS9EX4F
H7xnrdm5PkqAQwITcWtGqEPjOcRwXdPKgtlV04+5DOkKk9lu7hBhHlNxlhA6UeBSkzvqjDpcc9tW
Yhell9wpAikrWwk8bG2DdpYW9unh5Xveq9nph6Of0z6R+TD283AgQVC6n6PTJYvfB9NrSdP4BySX
8+JsSMCK165qhY8EjYz9mYfzeEpilJsdkX74lVy7gTQF+KSpf+ERsdbNMfEfyp0kVNvg6+gViLnu
5r/+IC1eyabxCnNp7AqVwMxaaWJaFEpWcGsjZiZVtxuUu9jLNnMxvcJkkY3GxwlliZHCdRGZTkn4
i3nF9e0xOGPoGWRl2N0PeQi0Va+tp9xrWy5D89SWlKI2k4sYiJPzTVVJ10uZwyBWaWVM6SSiURnW
GN03RMSkHzaZrZ1eUR2RtvEeKK7YAhd35Xpbf9YiPTy9KJXlBPg8+gsi6OhqbWj3L4Ll9svnP2XO
2cGbyZwI9zoi5LmBUbNorJE/JwHIKCPdpKwoqPAoJtAUWWS0G6zHxt+9VOhpr7cgsbW5xl4cBje6
1lP57vzVLR6j4UxEKrvOG/9AEkiLJg1nNfF44PrBNTSnoQjdUEkgn1qB00s2RmtfcF5P1/1BGUAx
zI2AH/OnGmFwefmyfL1mluLTlgDsErA22UrlM3d4UUL0nQRCODJIyEMqFzxZ41VcyCvZaQBHtP1Y
8uuIMDUBB7wzz6VnxPCfJNVWDytWBaPekgz5fmCoNfBIOiTDoWF4O+nL2IWmNP97cVekxnCysXWR
p9Lt8x+Y1ny5RXk/XF0waEngm8RUVhsmk3jMImkAcZZ9b1KHkY7o2RiWDeY96tSOt/ZXBjpddFkJ
RoA0v4qAz3ALVWQuOZm3dYDkWM8n4ZfAMnQwzH2ML3flwHQXl7AhYvwl4xCynofWHDDRehzMN8Y4
ohQipcA9fOgYSp1CoIuqmYQwbwE0l3U7eYIY5B/moaYyxhCJyNOQb3cogwqZhK9hgSfyb4eJryuD
7lB47OCOpv9Ab4ZCU3zsyWhzjupCut2qTqOCNUBp6hWbh9gmdDKMq7E8BcutAkz3CVa4tDDoj2dp
vlgDlBwEsY9UIlFDrX3txLULildDjK/LPXjesQFDzKR/t0WmWUWVyZHRa1nknDivjXyAO8LwFaW0
Umtxr+MlotBPsr7lIpdCiW7ehuzXb+3/mqEMWl8YP5ohlrs47SQLrd/nhwAu0GJXPKROixgrAlLO
WWP9bE/dbXsPOLZ2IxNxMWEd9u7HrHiLQhFQBQGDCUT8f41bRzb1ZE6LdT3jMGwx1pzOvD+jP0SY
CEEzvC/649lYvzex7q24c5BvLB6pO1KdL5pvTEktTaoMJifEq+6EfY5mj2bcyjvOrin5WGb+EPLP
3+6/x673ug09eSC2b/2oLdI5oYCr557z+/fFtTbISrurKgdxac2K++XGOzfGhJPERFtOw2s0KYej
JulHi5pvc8BFAmq+Y8HKc/cUkV5WCg+pbsqGvGXTp30fjvENFuKWGw3kKT69gIbRKgcs7POHIk8/
sMWuy045SPEv0sIjuH24RvQ1gvwIpFU0MYQkVklNRkxLtXzmJJTuQkdvW4cPZH+izIAXdMdA2M4T
PgFEAqmomunB2NOsAiC24ZB4j+m0O6/Hc1YUAlE7iJNbKEKZCX493gkDb5d1PDiHbngOhXdudcdL
jrroYMAPmUAUsMokZ1Chf/CVfbR3qtUEltUzVP8raO6hFlma74UVchBcaCcRv72K2q98CZkg1i8/
B6GfRlNDKOdN5t91jQiy15C3FFldoXFDG84hv6kUT0N0LCWgZHBP5PcvgBC37foV186j8aD+bjb3
O3mrsNYkzyWhX7nStoKO02kMytip7ofFzQ+Ge0N2uuLwloBBGffICCvCRxoiLmR7dLGtHlTzZDvA
bzSSH7h+dd6nD4jNy0+sTZqryqlPe6Q8gVomhWZicDWvJL9oj2BTaerTnm4HqYx6InbPBCuDP525
3UjYLybR0itERTqHUrXxRU/HIDJ0t060EXyswK6yqNQJwmKfTmBRW3BtU9Q1/4yRAdHcncAo4SFh
4u1smOL9JKUzTtI3+w+hX+B+NoEHuhhiJ5rN9Wj6UZ7Kbjd9nFvaXvR5CXJOXyqu8l60ac4xLiA3
wChLmhYVxCvP6o61M51JEMEoT/j3yuRs7+/sODriWu82Gb2BVgnwvgWiVFkOhoZawC3z51jvFzVG
+DieTmMsg+qClUuqx6LNNb0nJgvQoMrnFS1IN5witBqrvHXIZJKE1XlUwpPPndB24VMghE4GZFHn
Kmc9Hl0f4c5pZAm99NjkoQTwSwSE8cSC6rBZpfANRK9btrFvgbq11ZoPSvXBam4MT4N2v20c9FSQ
on+OQ7cWI31H0VqOaiFbXEcnFYbhizlbuM6deiVJhkVnhWrT68PZ+luVGO3ikvSmk7YfrVDOv3CL
kdRoJkR7Mjt4Jjdt4W7Vx8vHBUZmHJYdq7PlxmwDth3pO/7UH2+URL0yqU+Fud+IwnsoKJi4nlbK
zCddKdMVLDz0r47d8U6p+dilhUf/JpXLk0KpqiUFbZxr396AGaKc75dh6uV6rsyHZIamN2OWS1Ci
ACnQjsp1lGLfg86tb8emNeMm3VRgZsHl26E7pqoLme2jD2A+hlum/xsYPsn00v6oOpcracaD71+G
XNwnn8+PIsYGJGOjMeexPBlfJbsB0NrKNzjP9Ju4ynDjQ2CCCddUWHCRn6IWdem8gkY4xAmDaSHB
fLPBnOp6Tq67UwIUMp3c6o2bNrd6UHlvamU84wY6NcWPXvVNzamWOpKywtAUpy6B8vhpORvYaLAU
+lk3uig34u6PsN7OGYiYa2yxdWlZwcIrP9snAiFEW9lfZPmsjv1OTuECdBHopaL9kjuRFg55IbvU
EeOOlzgZy1huTRbTEchPHnJkt7wyCpWj8vl2py86bD84bkG6z+IjXCSCSvzCJMv7nLWgbjDJKe6u
TzMUJepj8ywRrShIprwSQlf9dQXztayd1PXdMXi/250ms7UE3d8+Q7n9IUq7p/3NL1+ImVlIuED9
u2qks7JVULg9kyAdN0a8N3ODPGnw5UCh4/dGQxjIThojYU9qeDWrd+ypQjpBodt37kZ5Rq66vDg/
X5jn9zSIXLZXgM3tSsO15fcA+Bedwm2doaEBALUX2P3A2S+CAQr4opYPY/kgKtTkJtUhR+EUmq6R
PG0DuThCVblNmITmmgRpxS1G/JwY21uJ89Yj0NV6ghfR99pl47ZtxMvAPIQODbdHjzJK1bWkixcW
bNhI4vuXeYSaLOCJTxDgaT/BSDT4JKzuC/giICnTZF8VCYTRKVpbXpeirOT6LjZQtlJxJI41PRHl
vWG1Ln32Gs+2y2lxV/PdiJItH9qTTQEpAaG0zxpuarTQpzFJ01V2icLUGQqyRW70bQsnSMBwPtNb
cbiatc3ZmsUWj/WKlQzZSjHWZftYTlXHAPAUCpTZ96hJYQ2Ig1by3l8AcClYHieGVs3maz93Rhpj
0xpJeG7KmRR3rKApEQDUDLAuQyRD26U5cs8Cp9an51MhcykjkZX/4bJVbd2Cqee9YZG4F+WQhU6z
iLkBIa7fl6fkQH6B91eSaYltsk30so1P/yXl025QR6NhoK1KL9c6+RnnUHHsVY2NPo18mStTcxHM
zirBCX3vUnkR/YTIXn1IoeXyPCnoB532+3REgsTFd6YSE7xu+JfKJ/cRzZlLEMpBPA6tyNh4lrM/
voxE5+0/iyUzAAMajiFS+gnuO7EAi1i9RB1l+bWjP6UwqQgzizrcAIjbiEeXxVGu4cOLO9BKXsvi
NXrLqLNjEXUpVzUF1d3ZNrjJcXxkLeHgim1d/+aeEjK5P9E35gyg+CHWvQx/NI44YQXEJygZFJkF
jHVHtRUuT15U6p1CzuT2lvr9/Pg8CZWD9jzNX4Zvlp9q4w7zBOnJaQrauRNmaTyC4W/pX4fcWVjt
Pb7QBb/lbD+fS2d3pUQqZHUR08pTQ43T5o+IoPOdBMUayYeleC1N23vDZ8cziOSP5OqjtDQXNKPP
ptaJcvurd8g4i1SPle9i8i4IKleISyPbcyekNtlD229PyKXNgwHPlmWI3Rl/+CGDj1TAHYv48nx9
Fq+rmhdjhW3+YyawCfgjvMFo5/+tC+a5EpEdfAhn6FxR28TskLtlOhZrq1eLDUjRReRRtllCBDx1
nFjAhW+lV8W7q4GlK8eFouLsYZlEXI8HbaDIjlE3VN3V0gmErnOzxlHJsBQ3H0Txz4RHyGEUz9+q
20df+elbWJzM0QAmiCsD07HjlX0SuJxxBTjHkFD/ipPfcgA6dLuPb0jclbaNESn90j1gXrSro10q
sQk8dP0Dap5VqrWTS04qrMM32a9NmRfEKMM6k1WsAvQYEJeGL9e2YiRK+VOVd+SXqNUR60Di5Jcs
G/pwirCkcnSQdy04TZX7erwSdUolYXWt6gPomungrRBJhleSrjKG/1T8gwMpx42S1nztxxFGYx88
lwdKYzdsbs7MQr9Wm+ZJhVdCcw8YCHFgeIwsd+s0r7i5Tk9mH/rG8sHLOpby2YEI3QvVBeJhoIsL
PU+w1+E/AXtix6VHWxPOxb30h3TfcsTIgF2N4R/oxD/W43M0TtCOGMUBn37UD8VeZeTUDXvmMv7f
OAOOP8dlbSKvUqzk6V/YD1cXnA4NuywQtn7363bHiMUtmPAGcwJuf//pjw3TvjWApLWzQP7cB/AH
m4E7ojAHCJbHPuNwhrLuplC5KSqi9qhnEZnMC27w+tspLG0l45Euvr5VqNdRC+zAH0e65kX07wT8
HgRp2KfQDRlmdLqonvu3dD//JiuBlrbLPWlMMc6mwgcJlvX+IEO29Bui3vQnlOwAHNvIygvygb0w
WT8ppRr1llozHMI9iiY8wzV/f/XT+VCLlu3WGeBCKmmIa8z1EYmERm7nnxFVYq1jr3vXzllnonSt
B0eWk0cz5W4BWqcnQysKyVOOk2S4ozTetXapBSrkNag5a08lH0DL1aLVKe1lSskmcTJPab+Ew8Aw
1dL9JyuFMJ8a3VYz2QY7a0BAcLgIS49F7M4pyRbB4F0tjIx+y3YDnBfcam6zqZQWMX5Tfgs88GP/
cMfH/9h9/r6EHNBkIc+Ln9ewvIpQEkERWSjPIWoD3B82MXOhLIYkLE6ykISqQEG8BvcM6WaK/i+2
5mKRcSjMWgiiIvM1D+hRgTLtRbJJB1PRPYRqjf7U/IS2fkSVZl0ZwHD1jq089cutVxIEU1CFV38V
3YHYfJKcJZb23RC6BSj2pjNlqOsBUamsEe4pMryZvkfuut40T1Fia89onNaUtjH9hk6y4lcw6mLv
zSk3Exj58F6HhU7T8H0CWj8KT2aCRyC8+3FOw53IDxk7soMq3eBigzXUtQhqJaKn2HlBWEyiT6aM
qSspypp95uP1esk0ZG7JlvL53gDP/Qo0J6bVv8kFsO9QB+K5fHF0S/G19JA8drR7Qk2MQfQJtiEc
VSHNFKoCrJHACtnFi8NxZaUWvwjW8ROonRPGp2XxoxVjP8EcdKJtNN+9HVORS/9Khmjpy3tf8eTt
o7TZQ8czJGsKpROxTzUMmgNK3V21LYavj68M4lwglIaTUcxGwJDGu4RY6sVIaJAox6VE9nSfIJFB
JVTl97YrWwR2K+wAmy8USmW0cd+rudN++FEGoR1fHoWSEtCQ6fGupwQtnm2ncZ0ah6bIXpCI1cNV
D8VHiwN8TOYl6glhfOhFKw+TaDO/m1xjJ1WOU4V3o320PaTluMkmnP3gVny900EOY2nsatw7R9NB
2no6Kj+JK1+W+4PFlJvrwTVV3CPn1oBXxxn7jiCsdZFMBKEtpJpaA/l5P4Q1oM8Ngk1XHRRjgErh
JA3/g252oDkqja2vJkgzzoZIew8uDNxQHPb/5Ko67jtIYqilMjeReKpKfDXAdwoEas0k2eB8czXt
jJrZB1IzNtGUv2TbXfe351JMR5lnrX8IUCxSA2BY/52VOFWaKvD5FUCFEoTQi1tB+juCelrjekzD
O6HdG3QjnG0hBgyZSWS+InRv7SUTZjroMQRWhcX+sEFW5ZZ5Oe/Cz+1e6EiiYHDUVBv1K/cBoyUg
ajk6+IhFUh+H3aFEphkh+LKhkq+ZLc6vRnt9UiWO4sBk7gF/AUr3K3uRW5YEf1pFVImMLGEGaKed
Lm2JDOHEI6J5Sbp0U9ceif0LJZLNV+2bi5gR4+ApjKOd2sijHtwcdZzAzgZAJTrun5Ic2lc4qqlD
otuYQxo5c/DGEwbQZkT47PGwpY7/w6KyimDkPwWQyXW4W3im4UCyX01EpgmovNkq+hC/yyT0BYTZ
ytYgi8h99ykGKD6j1uHwMiDBevQnUH9w0ZlwO/3vNPVOBfShyZXtwr/FkQG8HNMzrUfIY9WCEnrP
EI0imHb9uhQ2tMcN33Q8+5EIW7Lc5s5ow9xTABQXH614H9861/IIG0r0HO2yIo4ep6CGaKDG6ZJM
h979G+NfmknOOTQwvxw0LjBHwX/smxqEdFFLlw34qd6HDaHFKTazRf8Tn+b7w9WGu5gVcCcnJU5X
1GDaVvNxmX++936EPv76j+xeEzVCqiLOZfH0LwsulcLYdOxh+Af74SXquQUo1qchSRGvNT+ejDrm
rM6mGEq9vZsBFDFgV9IgjCeUvp/HOW1zUobCdPO0aSLKwZhPn8NxU7QtZqGCsECpdpo57vwIy9AQ
t5OMqptj4755WDRqat9BGQmLf7XQzNPXwzbedHXBYbgxCHNLCAxA3rgl6fCEFD3ZWS1AuKamXwsp
95xrhEBnLcHDdM57Zms+tmAUh4Op+wLzr5WCcMn5DxS6//dUoJdTVHvSX5ycmYC41502WnUCtheU
942W
`protect end_protected
