-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
U5BkC0AAtHMeviC1tn04JnKbg6sFZECbLKlG7BVI6jeTVA97A/EKLwlnWOQ6ICRLRcNN7heo7cmE
waewwIY2TNvVeIrCZUJHvFlUUpNVly1CWHqgX/w6j4IOnG0VCFwJiUJIjJ0GaI1rS7qLmG8QJWb2
Jdw08LT/PujZ/3bHsKyx6R805n5hBZZ16J8EXtwsMICyK/lmcd7WKGYCyNlSNfeuU2mxUMgl3R7S
0lh5T3S2SeiLcaJxEc6cuBrrSmJnoVvnCHvo7ukjGnQxsDwrNU+YzmVc6vfohZBzlkHidoGNJ2Im
YbSqKrnQW9xCraieVNDjj22CADoK0ZvPO3TQUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17616)
`protect data_block
XdroC44ejG6kAMhzaxYPJyLOlOFZnGO1lw86NDJLlUkAIiHZF8G1DrZHbfoNkR9138rHeU8zzN34
MvynZGhAkrWYuhFPzvtIKeMwAeAcb8nhER80eL7Pq5npYmKs/0bXDiYQ+YqA80BnbFhI7m4wyGpi
3QjJdzDK1q5kVJxKELuzBErGtXGAPLYABvreYbFZ16paq8SCUunJw0cst2FOW/GZxMXR9hgfFwDh
nJc9jkw9lVyt4692Gv9e7Qwl8XnCJxz1GkJNBk+IETjLgKkrfZJDF6Csw8huQ7eBFzhRvjnI5Bez
3BriCIr53IBGYGYpMq3EW/sAHg3FrLHNCI9Q/93MyzKo4SEw88NYh1aZA45aGICDQ5cDNmMp6fwI
aLoNxICB97eu+WGS88Ad88qGzk3PV8jl/jxcG0g5e1VlEGhQr+sZUr3R/UEQFz2XcKgYgIh1gMux
qDCd+DS1NFxplfaoO5id+ZtudhoKwGe3Rtl78WP00cCWs9sLaHT+hDzz95bxG7NGtlzWU/2O3pzy
7TPwAVBro5FZ7Afu0xmEjB19fJinAK3nZ6zkqVRCGB+1yAQFE7jAOlLj2su455z3kI4i8afnRO5X
nWpusIhJlnBAHJx5h+OKddViA5u+tFepkimKjfzwwR25rScD40GP+6/xiXLbSIPYhAqlboVZFEbh
92qKxJ1z5GLhi9GQe/dfr76KBicPo+ybL5DFN82HX0bTm0QR1A599eE3tdquaq9jwE6kVsGp9eH8
PL7iVMHtlMmlGxIGbm7XNFaiEgZrA++6HShSQGfFBEwMv8RietoYPD68pSkA8b0oHw9E64qHgwWi
tnClfbRDEVXD76AiC8IUpLBqdil1JBw0NiGs/d+0n7QuvFt4G54TX+7rIXCcQG/NlUx09vWCIQA1
Mfj4VMiXQcyiEpxPXHHy1DdOKCQz/lBEoO/WI8FzWeAl+QUtQsztxk0uiF/niI45UNd19r2yNPxc
ZdQTPR5uPn0QttXXpyZm92Dyo6SF3TmXkOhf6/F7XRt1qP8CznCdZE+6Wfj1MfIAsgw1cgAE/Vd4
tF8XbjvIPRTdfcxcSYdtxzanxpEo3RR6ynCUq4N/9PUtizJrF3zLar3XFmS/40B1GeO5fnp/Juvj
CVPRUZYFwsryu0AZkjPNjmak54yo7l2JrWtooWn3XoLuEcOMZGzLvInPchxQbxsgiJq6cEd/V1lF
rBT7Rd/sa9uB1G8POyNsYhj8HIROrrGssefE391BwgR1MqyvFrB6FWOADrxKgdqSKC2V//fae5iC
LSEyG0H41nP9bwRpqk1JxkJ1BHqZshLBGsmXEm+8JBcIy5xGn8SRlELbwHudY5G2VcQbcFUxN+Ev
e6vyk8v8bpwnOT55GulEAsiOyT8uZ5QtegdRpu6/+f1GFhfyjCtjUGfB8nXUQz41D85UYJN4bvrT
Dsk6BuJeIwMUA+pf6733/QAbdHmuEIk4WOgkiM73VoGevsWE+06ukSlHy7tl/f5sUK94JXTZFjK+
aVgket0bBHVq3QEfpB3z7JHa5xQkUCDAQzIQGsDdpqUWZ8ic59aZwq9nXMNWR25V0Uat17tNrhwK
PW3AE0Rdb7zmGpX0Fpni3BD/i20Z/XLgrXv+EIe/izMpqs/dXMs+Y3vGr0+37vxvV66ITcOGmaQU
QcKCNFA3CUT+QUBU1s6fUZGwjVp7MtuGMCGSfwNUZNvItDHaCE+iGT6aUV41rWQhPrWzIY2/MmqO
q2cLcis3jdR1JCuMStK1OVOYXhkBdPOYPTnQ5EhmRAhSRzkugRSf6zepzgbl5HF1pAuMDpNvpH6S
OPx6Y2qWZY8KXQRo9M36anLQ7xp6LIUn7ZL6vKwLebbP9CWU3gNVjVZF/h4ms/ZAP1t7DN84AwaR
Z8fJgh7YnhernQTwoQsjJmhdSjaqV8uxHhPW7KmQIE+WOj1C57Hwugka2MmX1zD0stnyrIStlesD
7Sa62EFYqyynJoSB9YOI0Y3GzzeX/HPq4XNBnMFsLBT1IWTIOPROrJsEMHc5Zdk98mZVfxJqI3tq
DtnyTCmMCnucoMIhy1F7lM/ZQ36Ro4P+zBsRGEVwo+27DuNWMWKPYjsDV3bakCQhw+h+tK4k6tMf
HMCwwxZaeBRbJ7NVRNPKm7e3Sz2LvTb80nCIb1zzqWOBrK2N1q7UtmI2tbMmCS/SWy0V3ijyMbB8
VSm14V9A5jl5eIN+TqwkY2llnWzwL8sk7nBhd90J0rJmmpjNdKRNSWhP/vosWQydv9M9gRZBfDWb
PGWqVC4P15w6+G4Bl2HyxAqdAbfkpIP7/dfNXynskpSRqL522C6++4XEHK+xNbfm2jNnpPDKVNr/
p/eVHYI2MqxVl2TNDZMYDgkkml5RkKpecOaKUtK1e3On8pXVqDY/IIufI07vRuYBSkvrERfITut0
r+Kyiso1JCeyMrSomsAihdmWXZcK6DjXKlrsrT8TCS45Mv+ctHOEPqcrTZEqNq+fGrrQKAIdKzsb
APUf3EzeyrmD0iX+L92XHx9ma6nY68AM48rgRM6cPevQOaoZhYuD5UQrCp638Ws3XBZ5Fuc/Acm8
j+er3E4P1elcyZ8CZ2lXkj/h0LvL1LmgWOHT+WgwLSsdVZ9xAU4kR3OjIh/v5YCwX0Xlj3nwLXSs
4JG28amen0pYTXCYTeG06h+QUgQB39IWu7bJq5HwnuBz1m/vTeQKtVVtbXooyUfxsxA+v7E+3ZRR
+f93mUKRsPH7jN7zu4JHep256UZlHhzru6saOYuao2+Fhk9fN4Jx5UtBHFf6d0UpKkRSnL/h+pcB
b7a73nCwBOkteZL5tmLEdykv8p2BYe91fv8LjvBAWow6nxMBX7jCL4C21+IBYijyDzWN/l7mCZ5c
GkuU6JAdnTR9Hgod55YDE2wMWQWoaMS7HmpANQPMR47dl4Ia/TJrB6faHfgWsTsUYLW7K6wuhlje
iiTXFY8sPpvw408DF5hZYFLOSIrTE3bm8xV1sgRG//P0zipwe7hPHFsEVRgX9RknzhuhIKX9tNa0
1SOtIaa4/j6gDvZ4ujmZmJS1GMkpgIAKQI+Ujh/gNeJyiYxYI8AVgkIOijwuPsE6nvNDC04HY+7m
CZrVdbhdgNgrcxqT6AdnfYn6gZAAJmY/HcgCSl6zk9B1A1BlTheODfYEP8Mcu0PXnj7I5vPCK/3m
80axcduNj+G8AKYjEag75idICJiJPTeB1VhbP5S8E+r0ptjSP1lNmQzm+k/V3NEMPc8E4x4GguB1
t2Iqauu00eTBni0Q7RaihajDXBeu5qTd04RAfZCX/fcKGWQs1P4qepxCeOmGiflo7qgKF4kWTda/
XOo84qXmWHgEdNuOqFL7Fp2V1c1S+JwuNAW+gBUr4pZqPTqww9YxVyfsrJuHIjiAYYAMSmCdQcBV
p3+DUdGPIn2n6eQThD4RG7J0dUzUXrx5xUa9WodzHweDw5tulZA5qPPJsgkcyU3MWqC+Jq/TN4ZQ
dTPrYhlKDtPy09dGirP+Vm6UeuoveevEhXNKyDoYl8noJWbKx+fcHGSzp0Mhuyra4iyc9f2xf7y9
MeqT8nKSNKh1xlj7vAKqAX87D/kYYKbxdIyDOPKDlfZZsA6AHm15V/1C7qkfdDHuMM+EK5DwcTNT
AYZUrsNARUrtxpgd8qiQtTHO/3DG0GOKbq8xtMMaikDoZ3T5DNsyu953DdYUD7XdtDV6FE9hcvpb
zsBmML1/kPb5oyhdTy5O9gR7V9O+QaDNAn7KrfyAT0MMxm9ldgNM5HZJLvqTE7L6cnk/zz1sIB5L
bfuk/ZL0UDogmASojW+4aHqRwZra3vzSu+RaWP+2EQO6eak1vcaz/WE3ikzVsI3UCFxlIp4dhVqD
rIAZSRvPY80NAl/Qf5W0JprqTn/TQkB4FaZRn/6JbHWkOyuCYIkV2hSx/CXNqvXUeq+tmP8LRKvb
UNu6zHe8IpqH+A1pB1QGLtwiBPssVb/rqdW3ZYhou60A6I/BbrXtcN71Ymi8/QanRUsSFgWYX9ne
Pfjlyispd8FJOJwdR8MC810UMMFDFVSQMvnpYKMHRDeTKP9UqcqYZs45wyfLvXY7n1UWp+Qi1iz0
mJ67+TP3zHB8y60QPapIYKIaxO0V9lRHubg0XxCMuMtxy1sqPrclTjmaUOia5EY6S+vCcI5duR0x
A/6Fj916L0YdqG9kvFdbKcgqdeXRcWEssLUiFgoXzJFY5vMP1uzi0Fi3bADMqj2zBWFRhNEixx2Z
EJpy/B9hbU1YuKg7jp71Tq1xNLUOF4NhYmer5wVDuFC1dfp0Dh1Vt+F17d600sj2kaKyQ5416a/E
ae3gWRKP/FymmG3k9tnR0eYDRsckWlmm9HF86PXEp2GULSk/+qodJ+OgY+8E3/3jT4cUVVtngWIV
oE4ADqzykiuWJrbEsxxGdNoIDMVMvh2h8D7ZkZOezyuYBuIb8rR95WYfTcdOLZ4kzC9xa0zhrE5I
YN97lUIhvasksqwclgBf7MegVUWnXU1p610H1lNy/rszwHwRoqevFsiAkLHJV0N0L5ZCy0g8KPDT
j4Uo9rK58HMfC5wXuVHZn4a/ABhBF3QVi3dgpmcpTGfe/ueJfKxHBHOE/+Ppv8/6y9OeU96o5Pyt
91X4zHPmQGf6QkHvhqfRMXNK/A3mjKAeA34oQWZEOYtnVqyq0be6/QURQLEelvJfih/9PllvvALW
ZHOs+R3iKTZiEAr8FMk68W7ps9OBbe/a35iPIZ41xCHL0fh8EB12hEH2yz3fGp9zp/DFYmg7hmYi
89rFOErIPgphKVJDY8wAq7+7IweMIArmfIfjdAJCyneHa69XmpbtQS+NwzcG8kf3N3IHMlnGpKqM
Ja/dVDni32kQiUnQNZAuDoovsF4hS90QOcwkgTOBOQg004pJerEh7jQlo6TQF+fgc4sExMifoCit
P9Ju9GHha4PR/VMSvPHJPVzUKpdKBaHhWwUXZlvTDRXka7MrvGHQ4zQHUbR3h8apEmT6Nn+Aaz2W
oCDBavPzUzXtREG2XW0r5YdP4eWFzsIzqk8i6g+CuzpbKbVATpVlC0GU0DmIuLrB2PQHdV1KS2Yn
yr72zJLZB/f1z4pCIGWBvhRoeRSC3n+poQ51AS15YdmAw9PCiHjINuv3aB5RfRvlCMJFp2wWle3U
rv8PpOpcccWWzilr8mPDjc+iQgEee/o4oeHg56F8HnWWKUKjpDAFWXRvtjzR9U0fAJ4vBYVRhPT1
fsmOm0OWnKuRAqw2jzpYvpTqonjR3lSRn21QhSFO0xCwDxugdLd2Vtg/fjhM04tLNLGs2z2qdsnt
RfdDWo7D4GmdPxzFHJ70+LzvjQ2aZXJnyjY18OROR10wWkAeeov+PHFVSWV49QR+BJcyE6G6Lhtw
QjZv9VeQbB/1TFsgv56pJjTj2WN1GPq4gpdHeEQrX2PXullagSzhWIOcQFlljURT8Eelculyls/q
+iPVUwUehtDu4IfpaZxC5mYwAdDueE3Ms2pNP4jRCDZto8KUEFIpDSzAvbXoO1ObZyfk3Z1ubm5O
4s2m8QcFcwCjpV/+QpfP927Z93eDFU1vqFlnIOx8rFRtfCC+g2KaMYAzQB07ON005qzBOCII5kvi
OaututIDHTiIRnJZc7zqvkGUQmvdCSElddbGJFn0vFzWjtsLNKuPGxO6cHzYDnJtkelOIREmnGu8
flumxO6zO424nV0qHBgmEEabY+54eRbkA7E907z7rAH+ec3fSaJdOMwxd6PHZXB0hlL/+3x5iEb9
JKedeBnayFFT4Zuc7KBOpAuPEhOn2jhpuDstxFt6IAM3rSD6ZtwP9B5w8HvPtvQ4bSUM3YMaM97R
O/YBBnl+OZc6JiwJYvzEyzdlfkDTce6zhNtK7UONkUZKFZWnHQOfIKC0A0HSvmJ5Wk4wr2AzBl+y
m4Ttborkr6LwXiTFD1wh08/TG7hknW42lQFzLATyZTCX2vq2mLdExavIVn8I7SpTeDzpk1V9/sN1
ibnXx27QtmIrwIcW7Zjhkd79wMaXV/PaTZZv9fJfjNO+g3kxjQOfVdGBA5Y/FurvOlzGD9P9N3Uv
jhL4SWsuuDGHexiUP7p0aP7nTDtvmTocRyWGRXkLZq+0GBWApdJ9YC7/LqWbUjHh6kS6t67UXBx3
ZXHPn7T08xmZDYQoZ+5uEpKVRamzo/H6yQblLfZyUECKg2Qd4Pjlkt46v4tqzgNAdhaz4pY9xJA3
MAEbZwd0lfZmYFftF/no9eq9G2i5qS3oQ289bXybwurAJViQBYb9vNHTULgKhH1m42ZNwz8Yfj8N
SdzOys52RhThrsYjTV2xeHOdQ14Xccxq/RIq/YZYSzjOsU5qBj1z8oZgFBdDP+AVUhmkNWbBMLtr
1D/kmFGFcWw4XWxCMb39+7DS8IjVWXe8r5BBaWW/bWAUwAfTDRZ7IZQbPT4LpM8xwKK+3DBlAiNQ
bmxdbyvBuydAV6whN1vYksNTCNN2ZnqJYnzCxtcbbPDaFS51jYBNXbEO3hLDiM0+7hXiD8RmHT4+
K3KTvqmIDV3q65o/Dw5Ie2urQz28vxMmqg26gTiSpI4zrm12VkicvG0aSJuHpWgwQgEY/Z9czOv5
FEBer/2KPH9axeT0u0ysn3LO16TErSQJae1Hns2UduiRopNlv0zqjeBIDJFIdv+do7gcV4pmDszj
cwrsjtWsC8Qc3sZwBCji6WU8Igqvs1uo+1hLKOBMR12zjQoRQEfBr3totDE2ed2CVK9bS84XMp5K
D9W6PHNmyjB9XIteFA4nEbVOeABSZDLamVqZXroc8uk/54+tenzegk5Ids4h3oqJegtkiGzjjmrS
Q+l7E6ikAze+otDEXvO0EM9gt74oFjHs9Dlza5F3XCAAFE8cxZDOHf+5kBDIYOHbcs4cj0RxJD42
2HKg82JOcdnpfKx02pMb8EhDTHsS7PUS/AxSBS3r/0QiazIwIaGH6S6vIZroAz7LFAr3WbdFXWvv
GMzty7aV8zwQuZNs1YmdFSarQa9T4i43FKo2wZq1O+x7iEQb4AWqbj5xruPymO1pMiMsgkO6YtHO
A2jNEXtKWXWQgV+C8aFaZg1c4HfT6oYIs7rTHXWirZiuRZedsy07RlFmJP6xuj9pcdp9OLzqtCg7
x783OJ7c++nT1ugqrmbgA1u+tCsSBZOa1LwKoknX0UI0BbSbrm76dtEaZ0AnhtZdEhx9F4+dWYQ9
K8x97L5tYgXNnVrqw7TYvkI+UQJpWa9JXdq33o1UtvSKYiAFdt5AtHYnTm31TDEIUSjqOI0uSggb
5X9/parGfujkdIynWXvVia07/1RXzil51LGaDL+QcigWbB6ArAK6a2lfm/U3QNyOCnBsXRWnAYsd
qqcH3edQrsa9mEHJ3vLYEMz34+Y5+Q/tXTsqRCKTzKTzVZytabZS7I8LcTjMpAgTt+cDPiURtpD5
V/5Mu41UF4likc4P4XGxmNPeiPrGstLwdCMrZ018u/yxi/KKGJM36iQourLYvoGKZ7ogN49y8l3A
+/NWgEoH8nDS9LIEzQsM8beMvfQK+TeQgan02jivFv0V2BJtlj0+cvjhewrFDOXekz+mOOBYpNSm
x0Rrmo859ngyLob7x20es9o8ghM6g7jYsZI4+3TT8TktlSA6VVftQzBV2CVBXK+F8CRGkrUdCOax
HEdmHBypvBnd6xfMW7ab1G3Rhv9i5vy/g2wR/+FG/7CTtZ7JBVBLCo64PxKvE/fzROAWjgtKdWOE
ClN9d8DhBb66mTAzq74M24fJmP9xSIM3rTWxjdhDflB47sdMDy2iOCLpaR3ftz0wVfjfPOX8aTwx
nUads1XOyzLe4U/MwLJ4FwDPcHrJnU1KTmn5cwl74p0Y0zwr02OjdyZIahAGg5Py0mbS/HIpgxBc
kSOFdUU9ZtlhQa01KDJ2+MEFTWACUTJBevo91OD/thsbgunc9RWCADHzThjnL3+ynVIoNqDU0RZr
ClOx1LvDQXsTmyAflTx5A1d0+SHdD9zFGhdxS6MHfa8WpL8DPZANv92+DXPEEzagXlggjKyOP3Bk
7w38HaeMIiVVJLXFBChYg7+ovHb6Zr6pZRAWcMNVDc4TCr7gEcgRPSmyXriwPIL5KgkQeaqFhYk4
1KwZFz3wcv3byVuzvMRaeK72eeglgkMJ2Ur5Ei0KNeaOBrY3TSrpcOeca8lfIg79cLjQk3hM7Lk1
NOkFIYscTTq1ajJgUiVKl2/fWmD7wSly3Nr6I0MoRJTGjQ6NOh8/Cy7Ft9NJhMu7SrqvU9wzSzpN
FHNTCrBnjXrQcn/OyJ4iuGwhM8UsZoTfCCrEJC52aa1XXR4Fh0V58De7cZkPIRtODKwtg/rQCCRR
BEPgIEBAgj8iffSRJCRjS0aO8tgEwnZNzZNC4hdHP4Hs6RoGM50MB/lWkJGDex6blPXfXsEUk+Lx
4Vbt+FQybnJivsYulwa7AZIMgiGn34oTCyFDnb3hr/mW24GqXRdCxzjPpABi69S3P/dk3yBvusis
E2b2M5fze/QBgkIfnhxIA6X2xoLf5hJEnP8bazNLZA7jdW3RhqS9QOi9//+93XNUw22Qrf5E24p1
1teYTh+EOo8IaPb0Ti5DOMDIDbVsBmZTHL4pcY+JFykjg3lxxD3lty53HaMqEcwpaMy4CPjGDH5X
JKXNE840T8tUkm8iLvjTJbfQg8EIu8EVHBe0LfTJGVc7OV9EvkziI/ROFFIgjsVOTGY7zPA2KNd8
FObc+Pf0ldZ4zUjo6hXOKyb4aG9l3dCxiqF96T9PW+bZo6ta414EmXty4BoHq1AFWqBeEDuP9FVy
tgxd8U4lc48ybaKqpbgpZc4Ob4yPpsD+Aao87eoOulq/VX2GLpHF5tETRh+pzAgtbr4bOeD4Q2wm
7Ua36I87ltGu9wPXF68teALbDoBl3dm+iF2K7ZlyVuZV6FMiUPbwfSrB3WkUnEATm4fkrskp8I7v
6t+vKQL+U87Lmxtwu1NobIzJT0dEWXZRuKbM5jW5auQapFb+IkjZDualdeozEmfgHkEXtIap0IkO
Q6ZwpdwEJBmXUBE6Rk7i2tTy0R7xXUKqWMwz/NZKWtQCCyKcV6oFCUAKpWX1Q7Qc+80ctq41UpEf
B1JOiZzCagDdu2L2PnXSKHsfMOzJ5LFv/AZXxK5l8TCDHBe7IWLvljjRXB2cikWR6m/5zLDDtX4b
EbTLHDETjp+RQA6QNAYoOQa3LcizPFSSrnE0aRXKeg7pRQA9eZKY3C9g4M6rJwNnudStCw8e++JI
bjXYGXF/TET3KCq9ffn20eUJt5UtG5wC2G4/dzmPPmmi3PEGzl3JcKZHNkqSfOROF4AzHi2ghkgl
zJboxlArGhv3hIt08tf8TAEDS3fP4p1DY+5P0Vke0SoQUEEus5Qw6l9ewOmuysYBgwz70i4pXkY4
XLbTjI0NOFnOPk8zpy9cOrMCzwBIMRbHMb09qOUx3zVOGy8Q5M7JtYUXVfedM9wwG7O7dRuQsTQF
LaRW7aEMTxFPFttZn9XkqXkvhrM+hYS9eYtzF3AIikPlPL0tOq8OkAkGAoPVVy1YF0+gab8Qvw9h
sipOvdNoxnGaYEYTBX4nSxtWnKnKUjSSyPS5EaqfHDVf8412u5rgQ4EyalwPtoVlyUDxP6vcBmx+
iGtWQSmXUg/j3WhqOeY1zGjCHfO4irM+cTc5UcyzmRYDukoeoj2OZrmlMthnvNrS1+wvAgcev4Rn
+svG0aylpEtHWLMOS90XIDMGLokPujoUd+UEHwinO9sTGNAE0TkqKzcYnNYUuD87uBKaqgj9PB8B
rrEwViMnL0UjC8zp7hsxZHKo5ZyBSXaSDVTFObyKio63jxtB0ClXgkII5F7EzH/hxkf6HgOZTc4y
i7S46IGAOalHNxh9K7q3d7fkEHyNHJqtugSlW3k7FDJBEQDRnZTY/3otznVGJ6nLhwRryWvOEKfJ
TKGydcfeFb9yLhrx72nf+Ny7G7D2FUqwm7KyNx+MBK4g0KbgfGURv89NBi8h+7gvmolXfvPTXIpa
P/yGB7a0IpLNNMi5NVOCBBNeiOblf1OfLTJNR4F3k37/6/hrLa87ahZWHPMDWt/fL5srBArNH/JS
/UAGYaygWdik64FpyzrSDMEEHIbLa9BQNmlI86OR2bJvhpL6v1CRV0es4euWfsW59iRSV1zt+YoU
psENf6oc/Qyr5teHhbW05NbWWofU4IX4BIbusu+gQri8vsCdxcL7JKbbJCAuvcg9oRo1IJGdvxga
BsbtKcVZba4suSxBJcrsrXm4YazY5gE0bYGfnGjYAXWX2xychKFglNt4gseTjKa/4qJHFbJ68Tss
fVcCsEZH3ecXoTxPDflHkGXH3/wRB1B8SHZXK52iTA7PlfcZ0AdamnZ3gwOG484fri3sH4Fxalyy
Hu8xRBWhHnXSjRPQB6QtCm2qyZLuPelz6HQmXLGuy6SJ8ceLrvuEst4tHj8NW23YVja8s1Pd5Rd/
arwPMlhUFoN3oGHjfyenjOjEpGjGc8/ne3yH6YcaFBlPRznW4OHMBNvYNUgYWrreMkSBDKsGBbOA
0Py9+0jNCzADwGixmWMS/SIae0mJ21Ri2sLIoAC9+4SxFUZbKEsppFx9N/e8Qed++tuCSz5lqOum
xL54vhENne2rH+ZdUm5wva/P2Hufymu3lOduxiWJo/ff8RBaFF+zIGrsrEulEFOZPI330sOrYnBB
laLSfKT+9YuJ4hj20GhiRYVSDwTWT90ygaAnqY2fkXDxV5mh9OuqxSPVb6qaqTDv1UbBO41HdiQF
1ClGyz9MoG10PExLM9hueKXdyyeD2uSsBrq/HcNVlBLIlShu9hRiCAV2ofuLAivLyJjDI+lX8jZt
TQlR4QFqs+H9Hkm6CuzKJDtiatwwb/KmLBnpOZCvRBLWOpwMEj6eSC59f/aakw7vJvxJQeOx75pO
9kGjMNwkRh5M1J66rF2M/XAUvUcoegwt/uR58C/ch6jZxnB/ddk+r2PtUPRGEBlbMZrIp12bxtXj
8kd8Ol1QJ+i7tkrcXAWtvBqztI5snWyEd6n/ecN2kf90PzQn7DOhM12BMgXj9J+p3PxR/qBd1xF3
NHGAi7KukXD5UnFZPoYxoApTJjWv+sCc/VKS7Mk0+UlFXcJjiwv1zveHuACvH5AKrQaM5cKfwaV/
g/2fzpApYIfj5QAdUvL6a2sNgRaDTFwreNuSRadLiDCzsmTQSGsFDVeNu6opfl/OTuQtNS8JCSge
gl/zYbFSb1G10af+r0hxOlAc0zemjnB/uuwRQqr9UsyZtcKh3VKU/lrBkIkwWNniGv+mTXhKIzeR
rrWExm1BbZ1Vh891lcNf9uKt3LoqbN0lEiAPBJpdBMWsEbsAljUsYojY8oBPcfIAE+9iYsi/ntWu
55caoWUFRE93M7o+Y0R494f5srKK2BJO0xXL2gdPUYhPYHFFoHDKS8pCin04EvN7TQwubnwzo+s6
Ca8OH4Kv0h4PaWXBWKhesU6diAZPmA4tenRBWk4sooGhJRTohhfG5WIO1Ij63dFK0ouliuQqyTHp
4lFwTrKZpRvb8vNzgmrX8i7+QXc7olRvbpTH0Sbjp6QZxFNU9t9QKh1LmN8q6ZVFONU/EulHTeGp
DzRqmhF9Bs8kPc9oETivQiadxTllwxvwRQtWID7okCnVxlFwpGEhTM+je/Amo1Jz+NFin35qUeV5
zTZQvTAAJbAWzCFV8ofEqVvIny0cXxA0gti3PIPoLQQ3Nj4oIa/VcV0qUeE7ZB7B2ShuWOmZRaQk
uwiS+ro2RkY6SbaXKLQxHAnk2WZ5069uikdsy5noEb8yfPcIki9TvOwEg7XHyvAfKe2ET48iGjQB
1lR42eGEFutc4Cse8MenKQ5ICi8PqGGQzQxud0UEPq4cCAdnzTinwd9aZ+rLEZHHCEZtcXX3QBmK
hNoH0A/e45xiC/KoT5n5IS+BbrWbxhDYPxutW2Fnrx8e9h4sHJslaRCpmXfAZR/Naq2lPb/tnc3V
WUjlhBiZ1FcppaRVqzFb6jRUPGYrXFOdzzP4iBYPsWQF4blWZMsAKNRAcCNUqr+NJoTOaSRe8Tk/
Q1ALLCTfPCCVgCqpaJlJjWN70WGaK8qs9iu6nsFun1WK3Zw4N2ZK2mLyHbHsQXnDlwfkbHBqf7aT
TMXpm7QFeFvzKXdsJeXcSRk3DFxe3whu1gjFYNzB+6ABSnudmvJyQLcbpYkK7+ip9wfISQmh7WDa
UOQL8m/r5tTLGTeggzDjvO0aoVZYjRvekclo4X19NniH/T1HhaU14IXl5q9wZC6mS6QC5uakUd4U
QzA8GkGxWnvO/TJpkwrWfrLMDgOM875wUmzReqFF32B7f7wIpIx5rHOfv4rTwYVcSGdlGMCN+j8Q
DReJvhzd+tojcC+FZLqCfSvpyHn42Yds8C1rxLcfo5yqOwLFqlIAdArGZP9dYng2zw69Ya2hOzaG
LryyLmbnUUEv8Ru+g/cXTVziM4clpifdw8D9BQaNwBbQxbLxtbcAcgC30wbv+4zZ2QThaR2y2jfD
lV9D/OWmzgtF2Qqyhl5V6JZVIEp/+Azg7UytyXM5YeTS2vZmDWAP5IkZ34Td47sHrV2+lsOLhnaQ
6tkg4aCjg3BiNbHodH2BJTSWiPYb7zRLC5uRBmLVfyz2WO2k+GGPw//PC6L1jlyRW9dw8wwr4f1T
T5tyjSu9aBo4abkh7v0w5Uo5Zyu4Ds+Mst5Pw5mW/ZYCtbBEL4DHrGifRJXDxPBzyGQsUIa9ecsi
geyjLsG0o3TAr/6KxE6+pSCX0peKktzlR/UUM+gkC35yccz6kZRjHZnlVHWeu8GRtjcMpWDJW6az
l7nJFhhHZ4Ri6jJHrS/nmeocFHYqxvr/CpBlhYkXiPVDW/R0NZyLqmmvD7FVfIrIvPfNktow44q7
8BPzYPvtpJCt4MYRtENZGHu8n7S6PXPedGlz3ZJEBaLIk3/LdOf/hnCYuOB4CJkv6Sa5p8hGXxql
3KZ7P/5K5oyBgHFWiqF7XiL8aBBj9ZZ7kryjxOBhpDBjmL4KEd7h84vUYEuMxBg4QhcCx249cQ8I
lFEKuu5ItGHouMJzUsb3ZuPxffRlGtJmb+G1eJpPwk3ja8Z5hqG/m76HrulcpfWHJGZG0IXgCnGT
0/8/zXWpEijnlRYgTqZwl3ljxNykiUmW3kcbotjbQbG2l4Hagn2B4Z7PJeDoDqkKmtja8a5ahtkV
kwOaDewYMHm6WA9aqtiO21ivHUsR/xv98m/sKzBhai3kcaQqEeQAdDLe2JxXqqz3zvQ1QiENXjyJ
F7MWEOBF2ZGShs243TjPt14j7o3cSNFOZJBSboG5vl1W4zvCzmI3kcS7JjS7kwUj09DOWZdbkW1+
ATb9xglopvqOS+gulgkvv8B+e9mCgasQlLZB7PqPgFKqqt82ON3RyX6TILBrkVC64rhM9v0FR4LI
xXpilMGTzWzCzShbzj23V0Y8wOE24pimnxGak4NUh5gFi06/F1o5SAqhkHshnlswotG6e5hkC4DS
9QQRBWWfKf5mPTBeIDWQ7r6VLX9H2fU99aMzgu5wrKYp3KEaFA8KppM5dYSi8FNJF8g0HHIuixbm
CQAAEZgQBqZ+7jn8wqjisfpRobs5LAoqoAZNF60ukMhtqrklD/XqqWhB/Q7RMTYRjU13Ce/ygz/6
LUcDnBE/ju6U4cFwMmLbYwirAlFWNe8G2ViN7DGAqXZEXpolMW9z7THYj4rvdDP2daPJYbgOtZay
0ld4fTeXLejViQb0x65fLHw7nKSY+A574YZvjUGUJw6WiHsRWkZxlNW06Dq377RJHG8hnPatjQst
52OA0O2JL0QbsqlZJe0MBulZR2fSA9VTo1FsCEpNWD/M5Ne7cYS/6J5EnnNHcaa+J+sBsJMULXxF
aHDRPGoth1EfxZBa/RyF5i1oL1XY6tR/48qv52ZPdEpp1QeKOIWhL2U2tbGSGrOQiqnzCZmdA+Z2
aAQwUv7E/CQqw6S6n3uo3t/ZKCOtGOYtZm91dM2duYSrNtWQ1mTQKuWoaP8f0h6/ODkNbEcN8F7N
TE2nMwMent/4EMetC5DQ0Okk3WeOEHXYWl5DMwYyXjLG5X+vLwkYzu/YLTA5p7a4MlKI7R384bY7
FHhOQ7rp17lAUrCXOq7ZxvqmNlkN3YAaYDwB3KVrknpHKdd+UyjNf4BsDq7uJu7VEQwg2SI1UlpL
ufow50MtENw7ZIfxlZi6Sgm3ObYU7Or4ACuJT7MF8Rdk16T1rLF9/ludTxCYr0CNh2y9NkRd4xbu
76vJdP9rG23SQ+Mx7Bo4nyhd6hjhj/3YTD9MzjraXheywm5iocNBexCX7FvrhRzFBZW6GVNvMuAc
dNNJqE0x7n47gqadulBoCEW+41zpR9or77L7ykE3rerLwjQaeX3tLouCj0oUIIj2t5MBufWsMWuP
80z6PvOKjt/Bpgq7TrHIWJ9jEo/HbnSGzPyTeX08e+FBjuNvPxXbNVys902JnlW4pgYhjREmL4cM
Exa/rN4jhmqc/9DTFCybBhHlN/Ai3Trz7Ygo6JP/6uMg8IZoT1LoSZHR2fBLuPIMrsxo+JFH+/bI
xlrBEoMqNu7ZQj1H6v4U1MLEA2wyZvPUA4uZ+Ugcuz5Lsrk7fan61yZW9KcvLklwvZJ/aOb++K3x
noniORBvivzNXkg3rElGrgDz4SwhzRYzk0uUvCANkNogbLQB/Kk3JO3L8k7inR6Gw9JVO/JG+VrM
saH2Ur8ZffXtHKAmJaBlznWBT+jMUFUXEpsPQDZ/mEAw2G6ZrJ1IWd0Hy0fkB1FvEzhDSjm6kBSn
4zxLls6h9XFzMRXcW+A17pRER/nehW9tFrFPWm62aaR7KVPkwe2S8QvjXRHEtd+6aVdS44D4PKPd
Bo1vaLVRAL7TcnvV1h5+eHS1Dlc1UTl6+hL4BntBoUQ5RujUj2FMA0VQIdAL62lBxQ+DB8VHW41d
CS7xgqGy5WO549VLtmkQJaganXSKrpN3qD3q0fV8fkVjiVTnstg/KQlPDF4rm1ew5wCetrActgDR
mv5u6E247TD7bQRYD8cptmLjQmUK2qHLevIjo1mh/9WDiKXFj97KQVMMjQmGRcCubmNhSKsG1H/l
rmk/4yJZ7U2sdIar51UxXjs3d2m0n6CrWbdlxOAiiharGWc7Gk1lEM+i5YgUPshPabOSzcrvePPi
b3Nr778cEKy/ZibH9viHNq+bn7yG9wP6KciVGobgQUgrxrgq4M/JAXsCAHHBucZIeNq8dQDOp2vM
gFAvqG1qS4nsvwj3MTm8fc23KvBUJJ4mzYt8mu6Os3J721FOPfFDZP+4mNYBJTmbeEZT0xTZygAp
5T1VlSS3+/nEKx3SyWf0PidM3zmFBvGC02LUpyH5tOCYmZ7dnN0SrPbUeZgsVf4duzv0kNnv5GXo
yG0YoNbN+iB4C3rJt50iHiGj/NeJn0mkVX0VaTeimUEQ8Pq+YuW8joX0xDZE2fJRJ2yTrtb7krWb
U5f1W/OSpesQCjdDecNTeQqUtEUjIHNHD46S7okNb8hcPrReT6psi42P0wtEO5gwzX1RK3mY8Hka
WeEuAiFepcokeAmX+2C8eBGIPKtkTGiGMnXZHbjb1YDVHr1C3CNin/ixUAtKIC53mqY020r7RyxP
Ybb5t3v5zeivH4MAL0LDC+GOZ7gL5GkSvus4hjVlzt4mzNO2SyW7phY72ly8/zNDs3pT9pTHiSJ8
/vdV/Yx0qEyvK/BB3VAfAZ6gHpbqoNpYvIvO0K/U2WEPe4uPhg6m+AEw/BDFNRzv5+J2MZgRLinC
05mLnxiGU5apAJsHKpjN4Xg2mNu2AIif89EHzseOxtkYF5MiJ12UY/ZkhY7whZhHBEY9dFYgosP5
0nWcnRBlunUiHr7SVuXeCnw4D0J7wfKH6hHIATP4Fr1o56EpHWqubwL66Tc/aINtxwOctXS8EGoc
kXbUfJcNG7IMwmFlxWl+R3oFtJVwYYO21Ye4sP0dpT71uvZ8KAlvM8idIPrSc/LDOREfvkqrqjoc
VxhrbMDOo+ksbYDytU0Wu3cLJf15BThSJYDAp0Z/cKYuBKYE4R3iT8+9IzR0IBj+VrIeL0sT3aaF
cm6/vu+3JyT6QHiEAdWDOJuEaDH1JHM6xeLJpeeRuAceoKttUn+fCK2s2AV1Lnrdhtb62+frhxO2
tFJwt45Ru1ktXr+QzY42l+2Izn6PWd9oa9LELqmSUsYecPL9S2VlEvTEknYO5SkfQ8d9o4cppvg5
aAY2/68wQWybzwfo8jeWwL18z/PgScXZzXRE9D3TrTPTBHLwCbcoAjFdShJ1Z6Nc+RADVjTPC7+R
Ll53ILr7C2E6iMwT+EbnO+fXzLVj+UzCD0bRHTnSTunBfZW4ttdvq+E39kNCaEudtxlTiqZCIUtB
qCQJ6cAp8nwH/84/fW9er6k4OzbFB90AwNPnOIxOUvRQDjVU6KfNRQ1AoFgCJsMT3Yh0Xvd0nuww
IWKR7AymYv957GAoUcMQvTdVWWbF3BxfW/OoJfLJwQyJlXxtGYZgAS1xIHAdTzteJYgI3nNqkz7e
4Yh1djibXZ2bJ/XMfCllBHLCrWv6nYxQjxOM0dCA3CTIatEdBnB+7J1f3fsIu03g2M91I6O1DMcv
F2/JVx6LOXCKMyJeH2Q1wDRg2QVtl1HjaM/lkaSIrlJG0lujLevuq6ZhUZcAWM96WoqTWlEI83+K
NlmrTJUveFsMj7Tiak4yHyJMRfiQaanK25mxuqbirqegX8nBoJmI52AqTd4s+LEbkzQ8J92R3r4R
vxcJvyvgpqcAzbORFiPKV+TpHldtbLC3ep8pKsARDIsxgqp7DHkHY6b7Y1b+k/f2XONPWe9wSAQA
L8BO4dC36pwvOaN9Fwc1gDDjT3mb7FJZZXIY/zxfj7xEO80duZqUtgnct5V9Zw5KKUBlBNU3Wfr/
2LMYNApJ9qP9fbKCBNFkcpRVs23P/w1N0Pt37DZo6jV4YQaOF6LtrOMMjw6xkB3tP1q7knuLw7wy
tQ1GmkHGRVTJLjH2Jnr/kTr7YeYOJ7XxWRUYgvrjR2pqqzxi+mxUXExXDREkMO/Sc5Ss1KZY47iO
Ng1e3PRnryxUWEvcnTHVNdDWDqN03gyTMe2kHBL/Uvr8ppWAckEjaZIjRh6XlStq5N/5+zanW6dy
sC2ZjLjE6TBmsWML2YQL0Z/OQye248jwBnE6Vgl8KztGGKG2YJlkt+Zwx251AaMLiJJz7T44Im6o
CzHS3Yv8le4fgdR9HHMVb5lIKB95CKg7iMWK4ik7QSGk6Cg1PovNrO4H8pCXj2wvJIXxS9NUJhpp
yzsY4XGhrZWaKQ6VcwgfWjvrYsvVBZpi3p5Bq9odTk73dJxXKxcBtqG4NSUO1OQdFEX7bp/IHZ+3
ys2azwRolu1CK7H+IfExUXtSM0Zyz7tCqP3oiYh2GPCpbKLGzKYm8Yd1HjgPu/zCo54y2np22i0m
KaeSuOcjp6uOfSty5b59n1ICKZbk6HNmDA14rEXiUTybtHHQnx51yalO186/aM/4KWAA/ipHcwMz
2W7hlr8crxlNieLb1yCqmQMnnW5NHmmvW8tzO14t9n+Kjan4cLBSV6gwM/I1P7/Llvs4+OVKoLzV
gdXn9hP1+T6gHj0aAyUYFzuZZkRGJo0P6q8vlQxaRISa9uFegQC62c5RkSWzg5lU7H8upZOkgbDa
JJyKHrLTVtX1+5lo90TMUj9aELrVNMRF92fQ4GCw1q5FGGjg1fBS8m9hPkrjdItDbqcyLvOHpCI0
V/xrIoNCA/L1nCnVpljYg9uiqv29D30ei5OVO8UXT2Y5ywWmc6Q9OqZQLUuIqADiGu2VqA6EkZQ/
lH1YyOFUJcu+hWeROOewqisoJhb37C3xgFE6rmgH7F8J4gLkj12Sx0vhmCFy1lmEFtiaEdUFGvQv
cUCTMOM4zqW0lD7D+7pKHwHddAqsyxfJqvsyFQ6mByqGE2exmbZ7Xa71VsUQ0Vs6OfRQIR003LMu
4QCHoOzwV6c2O8UCkVDL/WuAzVE3228oGaWHshri+IW1IFWvX3mwH5m8gevX89jNetgczQReKN/M
yDJ/wOIBlNPqyISmmbo8BcsQAiQz+EMF1+GwnJ+7GCc0SLgSb2PN/4F2l4Hu6rvXJoPK0ZmK5ULR
Br8/gkiSyVgY3bUW0pFkYIci4PjWrQEDUJmhxxyAWbFYbQSNQ7qLVXS406OHw9MOZw0FiVVPi3ia
kkXf1iA+UzQ19wbxaNdmipeUHm0r65xN7Z173H6bnwOpHj2gEnTedAQrY2wakDU6O4ylqpfN1ocC
N2oxV/Kiu5Qnd/cDwCWCEBMcrSn9tJ9bVNFoi021KrX2tY1wZ3T26WpuDDUHFMYu4Ky/0liVHyj5
S1PRFhMRzstMLomYMNDbOWPY14e9T/dD7ewG4f6TJyp55y9ZHMiG1OUiPcs4kqhTQAGnCZ3rU026
797oUoEocbGrGahUIxhqoP5DWXsMImJJxxiJVS9LEDusg97ssVuXk8JT3M1WcmQk9MFy/CKUXQDg
2bdFLUpwCMhktClr9LdLv9VA/uQ03dbQP94LTmpvJiMBHuWXDZKuV8RvRjFYwKO8JD4vwECSKhL0
CH+lcIlaJ6p5Y29tf6FH1TwBtf9o42n6pSLYlB2coliUMiOSoPyoO2pX2DzYZ6qye1GJayVRpYZI
1EYf9T2wYx4MMiElDkdYxnXLph9KBC14LWYfpQmK1O/PGVpyiakbc7jUjobYHUu5fvNCdWqZCOkY
JzafZUG0WlNywzpYv+rnkTo+jP50bJ+m710uhZ3Yhavm4CxuTmWex7Cl/4ZXi9D9sspJ3o8JxD82
cz/8TMzeQhfDDMo47OBaHl5vy/7teCcaCV1hWF5KDRypsMoRyFrIjC95f7ByyHBB/6Z4ID4XIy+X
pkkLq8UgGdPvmoRwH7sWWWWzkU+bbDGNzP9kwzguOhsWINatCP0zVYDDx5Sjz9/l4oRvBMMQLKGf
Vd/Glpn6kWfH8rkzqiDmC+ycpaskvryB+snU6k8P8q0fIU098GwvQtmAdOcEogDm4Dvip1EqvYgV
fZgj1e27POWdK/UYoAeL71cRF3w6v+8QPfNiQxEpn8IxqDGXmh0wJd6i3Tacmk3HxHTyx0B2yjgd
IF6lQ9IIrZ3qcaFY8EGg8UjSwIAgta3U9vxlgnh3ItVuGk8jt8fkn1CN5RlLrpqzmh34Qz75igI5
EzQsWxrUwb5ayeTFXwFuYEEYbEpaY/hmpThrbMF0zzr0i3Wwj3x63SSrvn4pV/g5yOq7i7pO2krc
cPAPw6GJlTYzHZfnvWHKFcPbeTVz2wrjySr4qHxPTOT5hn4Ltlh+7sXjpDfdd3xRf/pmNzDrY9+8
Iw1s9lnMVQyEdCe5N8g37tPDF/twIK1LebZU3Lzj1/wBpVHZHiFvTD7bzj3QLGAdZ8YXYOxTccLi
6jdaG6ceOvVsJnYj21pptAJOWNrdfOeudIUvcapO0nT9HODnFYG9vsFrN1flJbEWCrZHoTzqWPei
XaeDAEfILhZn61apX6FC3xgV18j8tEliOGUCRf9HtnV0VC9b7AK6kB87Rv4/t4XHVeruVD7q5x70
pB07KhQUjkHhhOslfInm6c8U7s/EpKrd5CZk2QugwkyE4WDKFwPVPubCsJapkC0ng5kdsSE+0jqy
NX5nbu4l1VT7Aoxjkann5stgdn8xLLExrnvaN0r9OCEqp2VtFpeWA9NzrrCbwnm/y4OYRqSzxpZw
mTqfJl92sAPn2Q4zTKcbPvztazP3iumP4h36QsEUerQ4eRPdy4F/NN+J1dzpIDO9geH6MjlPllWv
aiL031WKTD3P83dAJY163LCujkwfAugYnPtrr0axDXZJPDzDa8qrMe/zy2PKnogylvJTULI3JnsW
iJJp62kGD86xU6JrNHvhpokjRzrOXhQq39278nObQD/lhDAKdymSmDP1eC+gIUAmj7g+lxCAYHto
sT25PoIEGsqOHYLKnhufjyN/KSWf3y7fyEXiXavvFUX465BotIyQzqMfX+0axl/IdPHbmyhl6zCo
VUX5t/b66V/Qa9p4xE773h2gfNpgOkkplxo1YDXY0u0ULiivnqRU0nYeQbBWDkOnxQkirpRvdLVg
vz3Sy43qrhEkxrhh7RdVayScetB03gwOfbACwwO6IvS2Ns0Dc5aqh8hnOG9SugS0Y/VEWAiiUSMj
VvzJKkTmQa6WVa8LOR8UaDPVxwFHERc3abeUF/2BDuw0ipEIHIRUxH3Qk5iarsiLsThXnOaJlryx
wZPGZ/j+/cDgVQZjaEi1aIXwN1AE9Qym86g8T/Oj0lQa48wVBwsgbSnZid9roTMxsIPn26KRjiSd
oMOxo7iI3XUctKfMqH485i9PHFgui8mSMLneJzp8p8GtV7FIhBagI/UZW61nIkX7UKLcWjS2nggG
xi06AKENXNuLTNX9LnuVpe97mTNULpJDGk2SAYHpjsW2sEAKzqYuYYIwn1nceRPDAjxllJRuOkF7
CvuQqi3kacqfxNLpDD9PJZGgNedYmJoza4kuCfjrwQ+PNFPygkIz50wYotmGmB7tfUJhCSRF/D/F
Zcy/VEA/1EoADDXmFitT/edsFehrfhbObi0JXo/CPdYK03zmoinj/jIw2tmMIgHyfU2my6G8eo2P
Y/lbumLGrLm1W8s3I3E0VMAt2W8P65odHoumGpFBL91x6MaAz0xKm+knjTRswZo7wHr2jTANBais
S58zBsqXsG8+wfgP2ISjJ0Ckhz+s1b/FLL/YwpHY0X3NQAiV/KotHWAZXg90WUAz1fHCPnQXxAta
Hl58Pq14JPnrKA8LaYOuqHlsJmC6PCfT1JfM0eZ+qjLeJDwCdpvKosiO79Nya03wcrxddTsUPyNL
CwLH8zzO9bJQ/PI8D0DhK4Fslj8rwKcPW8yqPEanp3BM73Oi7PpXz72Iljj6lvqTD3S5JFH3xxAE
g3CUgNLtYhGy5zg5Apc1uVpU/0UytV+1GghzkAsfqmi31GoOpagpdynGKAEwoAezxhj9F7iBJDvw
4u25wDG+J1Dh30SEMMYb3vdfmDqyCoP3KC6V89gyxcR1BT09oOm03miKvYtsgxQ24J2cnITPWzGE
ttbF/7+aXNTRrm5kFksuz00xY8iVmv9XQzQg9jcTg60RUHyACfVNF/tR1YxHbvKKTcuN85AmNkbh
zzSgJAh45sGzir1OCyUj9W0wlwgC2lFq6ip85mJJXkGTsvkrUr60OGPTbr3Hlb02nOXKCU+9C810
sfZF9Vfuisn1NZlD4XumlhsnQPwNaXaM75IxgC1khKlJXZC0EJ6cNkrzr0waC+sMXyQHO8PGwuKq
Vg6icn2L0k7IhTLHEACqYY53T8/h/3/6F2xVKOL+1bKIw4AhytdDUpCRA9Y+lihjB7GlKIADUvIr
B2PkdaLtbdPp6nDucH+xN3b1j5US3KX+uX1gR2ksfMZqhk9FbcOIfSlMk6QQ2438zBzR8iVJ6j6R
dIgMPzemiOiKrOEY8hIuQBE6UerfMU83pvEG0X4DC88cSWXEd+kSfPeKRrrGBFT1m0hA2iEQaRDr
HJkAALelmkfvUnG5wmZRjkYlKp4c5AlqLvEFdUyX2fwzZ1GinsNdfYy2Iy8/8fBGntXxZI0gjsAw
jkNGphPWlMOSNuxq9ijO2AxXgxE3l/bJpxVD6yonStLWJYfqEGP2tDUZWTEEHiFFGe1rLd3NlIgF
oLqXUicGu2eYCFibnsmLK0YSWw5DZjb+fDnbpT0nMPhB6FhSX2teOgTxNIXhjXCc1ag86rTLGPyd
SlhtPd4imTW2Eup8gvIqJ9u2yxQngq2fUgfIrKFxU4LQ575J/wJbXNNrIoqC8LrwHcpzM70aI+mm
DVCD7vBcGG0Y8R2m0R7YRMapY54pHDnY2t6uhiXsl242aiwKBrIIp9gj6Wu5NpmFVDA+mmN4kHn1
eDdEPzof/Jy+Py3rz0krH8WR/Rd6+rAdgumwwRuyxLu3ifj/HG31Etfv9hkwnJ8Zl/o1LReKyjk+
m/IasF5SDBEJLYdP0YeBJzFhoDibKWpTDnobMqV3qV1qq+LgvZ5flCEvGAff2GeZITKfQ3AqN3vo
GLYmHgAbN4qiu/GGgNtVYIbAhiMas/loHxYNQdc3Mt5+3qyOF+0amAtydkaKaEFebSwY9XjRLbz7
oimMRMjR+1OILsuWc9/+Dmhr18P3/kwFrJjZwmkQd12YGZSyZ6q96Ek1yTmS2ygBP7sO5ePXzHCN
wWjFxU7RzsoWnrCNGArwIUE/Bw7MnnyBXb4SUUtCEIUCukv3DZd2ZTRQGngpzWI+fqpyhNxl9qYW
Iii62qqT9NjlUo4xgWf4mDKI24WKG1NjZamFV/w/df3Y21ZsY7ekTTwSaeDUve7iP0zKLJHv9C0I
+qk489sH7m4IAx5bakkxFy4FcguGlzPmNcFhlTYF9VljjqpO92x4kJLHCSmJV1r0sc9GTcz3MjjT
rsNijov/vXWlI/Cz/3dDcKl5HkBC0oc0O4FKUzcSKR3DHu12SDV+u17trTBL+IlXnmABI2DVPIC+
1aDHtvke7c3G41eJyM14jYVFgAYZ+QMf+5e7SCrm69NJtGUx/Yv2JY8hN+W8hVqN6/AaZEj0PK03
nyiU/Yc4R4JRNNYmLx4oCs3Td6MCWNBxya1CEd2skdaMeTAB4uns7O7VsHhGiYIKrF8dmMvWxPeV
9oB1K6kWG8b1XZGA24KrYD1be6ZjPUulntDZPvlUqdyuDKCPPFZ0UUk94/YASDkmRNy7/u5+RDBc
LG7Ex6JMg63krgqCutaQNjU05nWLk/Ouu9TxOxsCHftk0kciTUVfRJG4/oPs+4ySgjm5XcJpSz+d
xhyrMk06llJimTVCdOA1XL+nRVqrWLD6Rlqw+LkyJw1uOAn9j6b7kbVfz0OfVInkPxRH1DSppY7u
Y85o6TpInhPiyo2oonfMtlA5fsNb5Nihp19n5AovHbGyFeKdmCnuyUFMa+Orsg/Bcsc3zmhNenEN
vDyPGYgFKrgzf+QyU6JVBRBbM6zsFuMv7scchNH7FnQCxmfKApmTmfQQa6RU9ITVhlkUN/9E2GzX
olOWmcTxDE665EeTR0YozPMpA4Pmt3Bu49Z11fPGcOQ4F2ViNg9zxQ2gZIfHDuR2fqt4a4a6kVzx
Uim9HJnQTrTe4Rc8c5VrMCiaGXIRpefu9ZkyujBNJDbGlD610j9RFxTT32bwHN2GOCpGjw8rHFdz
dtT1lciZnNc2CIX3Q+Qi2alhaPiSvpze/S9hyHMNWGBWGo7yd0qKv/bhCzINYqfh+3xqE7546TG2
mImdKrKQt0orNWniTW6HQsivGjyAGwdFP86qllJW/7Ky2TrSsS0XEoqa47wpG/aiv09B9PZnrFJp
XMTvcaczGVZbPozM06gOy7H9Sgeu7NscLHVY/awawWHHe3ae2N8d4hG7ijNkhiQZm3kNMPNwvdUo
R5T8
`protect end_protected
