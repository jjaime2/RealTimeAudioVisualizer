-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mAPmRTOAPLFTYgXMMgCrhOOoNJRaYVUBaazn4Z8ih9ygeM7eVbN8o6xCl2tRtRvs7+iZwwUHM3nB
w8/tyCqd1Izz6CgFtILNIdmlvumCwFmytDgqp8fd+jhUzNfPMP/sz8i/aj6dxzXVqn8hS+HE8yDk
wX0KINN4jBaaT3FpK7ZXl4NLeOhfqZgXd3m48jDENHgfyQvkwbCDH8bjeWJ5uJxf5YwVAkCuQsKR
EBqvV/Up6IOGiCitQ+N5mrp+SnaYIUdN83nOCjNKGlVWNauk7ROcVFS1NVAlhvD1KpJS95ui4qhs
mHZEBd6IEy3WevgOp1Ea86y5HYH/GHpAq7ZLSw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30816)
`protect data_block
bSHC8EInDr/u0cNjWevgIjpskzMbjB7TNenDAZLnCAwEjs4+SvWtoiPR/rlJKt+0X/rUEzkh8kPp
JbjhPBfYmS8DVLOhLGVs5ZzKPsvnE3pBpi+df8JDNtwJCrzXgW7YuZAEW09CpigeEPqWZ+1l1UVZ
lkix2FV9uDvcKQSSPIm9brrk9a/MX25C4BGq6eE4z/PVyTu5lfC42sUMy5r9NbrkqybUaYmPD16B
92aswS7eX8mN2tBdm4HuMXS7kqK2vn8rHMdyUJ5eDiS0QF1ZgTRB1yoMc+Ijui2nlybDY3l/hCfO
UohX5BHoM8+6ovm8kwnKDIJgRvlqQG54WdsSTxFUZy6qsNbaicIevwWQ0QMKVhEgokSZ5KhcLrg8
AzB4faCA4/bUfUbInhYmtIez4OYkjdJdeurxru+2nEa81KHN8n3u7LOGRBNfg5/ylyZmRrOKbz4Q
if6k3Tm1xFSEXYnmYyktWo5xjfL+tXaopzPsyem0HBQDd/cEJsaELGtky3HsKLA17qCfoeU0RGK+
Z8RF3+0sNAhDpYk5goQxB3ycDJov0eOhh3q1UkeT0wHqEsy8MeqLgjiKEA2BP/aMkEDw1fCuYB5i
YMq83dqRaFitqbQB8j33hqpK37xLwVqXJUcrdpK+R40cXtplILKsrX/ap9dHoHpQDDxIlgIG9Xyk
CrysA4112jfec/JjoZftaaYrelM8Vz3BhuwMiKoD0RVryOpNot3OufJ6wHcaWET/eE6M9UN2SrpY
9jYf81ZaZQ/Ibu9R+Ac4qtoq8FEgglZ8lkpQJTOWpAPdyNFa0XyGazxj71DFVyjvEcW8Wv+lOLuo
A2Oxlbs9kVEIX2eVhC+lA4bzSI91l4Zmwl2DoC83Cku953H8/amRhk6fh8mL6rG7C0V/cAEGZVt7
YE+1IHCudYZ075pXeFm1mK0mmyFHxmDCFWrfOrxGJVXq6FQpkAFWUYUbd5tx3HOjULMaCPQ/UDZk
wKoUr6BzoyHycRfnNMDv48lecKzztXUdgqyKSQV5Jtk4J7Ee/tt4DOLaLlBCYc6lfJD8xEukIYn0
DHpb0xzlEv5xMhL4XtUBjnNtkd76iisMlKW3fpajF2YmBN2KIA49J8E9oWop1HoiC65U3vpEi9p1
YFIgMx/0T6BTwPDn28UxqVmC4XQzX4HBAebNIKjP/b2Hn0gW8KhDRO2Kyb2GQcqxGcD6VuvV5Gct
UF5k+toSXV4m2MRQbGmD0PRIVcnFq7GRoLMdd+KSRLcrrG6KcXmG89msXVgJvX7DjRTZyNWi4Qa3
Qk9ItgkwXy9CiQiGRQy+dc7g+qHyfMMp/sW0vZzi09+n9XrONtEBx4mmCZOFvY6Jm2jm1qjpLgX2
XuwFrZqRRwg4Ok8fMgrw0vYv9YkDjW3WARvhlwS16s8/n9FMfgkpioOvDlS65E2rDEk1m/jlBHIZ
WsnX2wixbdwPTH4l3AjTjBrxySIpKMgI/UQBrX+l45dHnHQUijWD2jbNxUP6V+ZW5S83sZY3vRr6
KYyBjsuA6VA2I75mMEB8aOFkEOtL4KDM7YD1v24Gjnnv46eN4FsdsG22Ncs3XTGZwa12FItJ67x0
1UrPqd1kFsxcqJ0gd9XeBPeSlSLfaI7l0QHdgouRq+/3VrQi4zJdrTzWZTMXiyvKJsBuBaU2hrRs
fO7phJTQXRS516mdwhIYpwZEvaU5cvvdofBYBnBPZziNLlMZsJtDCmmXgtespuBEFyuZCjTcM5aR
sf65KSqo7dL5UZ5yTJzLti+o4YnM7xSJUgEMKZngBtVYCJTv6kqGGacxOQB0BwqmpmCloTf3l2mA
PX50qItFl2JD1AfLaQfi8/ufgqtGPsWK7C84/Lou1a2Rg8wT/CSqayvjbqRO8C1FstF+q4J+CGc3
MZmTYekzvTufWp2Dmar7gbfeqy4vXxe/XGH4xpDMvcPA8hZjqEs2Eru5PvCdS0fWfN/GW7pv/yri
qvpW84dWK1QLEqvkj80YVse6Yu5wzp7C9tmp2OzMAYxNxndGBndYzAvIkuYt3Ff2c/pizvm6TsN1
eskzfry8FaVrOCYu8TjCJgWMTB1mPw6wKnQgIT9qdT/89N4e9yECFbVrpfLfnpB3B5zJ2CzQw8Mu
KkjREdHgQHQBV1F0CVhYbEqaGHnHUuge/UBVzIAkb+dO46RFiNmVAVjOH3l8dF4NDvMUeSqISjd5
j82j55tj4eNdeVxV0JuNbpWQG7C+SmagYfb0wDzeNAcelyJlO6G7kxSOdXXulmFenm3sx2xS6K9r
eoxTcTZ0OpY1LIIb2Ydjq0sBgSHXjgrLvwPiaRRFcablag8bwDxYtTJJrGinSV1LN542gqpBL4b1
SMWD8sKHb4Ynn05lLqbgd9R2wDUafB3Zk4TCt5kgjChAs2rA0wPwzNHTJI+AxKmXosNuPy1jBxi8
c7UEh2GRV/hKvKFoYGxEhbEt4QLtPU1XKZ8CgoI25paKcT4/tuGgrMMjYwFbS1t9rKAb8EsZpS4J
V4j2E427XmUYqQneV5DLMgFxxSXWZwtKFxMSBp9IJolFUVp8JpyZv9zz+ygKXntxewXoYi2mlCms
chN1M1En9phxN+eto5FjgedTQ6YlqgnXVF5d+XGI68r6b2051vs/UcigX7EVsxxvf+lzY9WChgE7
U+R0MvZV4jZJmmJCRUHZTFS0l3TXQP4kegwME9R0IjcjmYauOVVzbVQ1op83/8RyVnzaTVHnVyo/
YumeqY40tiDl30e7OU9HCEdww1637+S6TjfV7aNuu+aPXbxRTxS1VrqX/yF4lNS5r55/nGbybQ8J
L6dAi5BJMEd122lRZcPTp4djxSMMGk/n/a7I0hL+X5ZZAewDVAYRlN0fp3PcZ2s+Y9LpQOpYN7Vm
zH109fehXpLBUB1VVLo3JATqCJ7N7TQBA75Y8Bi/x6xweQLRzY6PlNwHPJ468lQ3Vy6LjoqJR0Td
iEiwljT5xX6wJ2jTtKvhkLwKOPgVh40ctyvR+AsKtfJV/DLfRTFUMk0XFcGUbyF7sVgaW7C2AMAO
4y/YXkONdl6ZwxxVy41apceWNeQ6vhL5djkj/3516xniBj+X2tVUUcLD8cAj4yxnu96zpR8iscET
hIkg09Z8GtNAOg1s7x3gAbPIVLPnHl0QT4ehbIvnWS8KrVLdQHPta9Duadiveqw16cvuMAaWbAZz
VEy6osO1+Cpn63F+v2k2jv+R84TyYBDFvsip8ful9FN9sgWYZOZoC7xyrQ1zphBhoP+cn5rLnUlc
kRQQq2v4urJgDBmhesZR836c5gQQG/UIRaL4KpBJW0oCNuEs83tJtJQfa0elbYopHFmvXBu1bcBP
jD5DM1cIVjTVbmghgaA/IAsh8FzsBBHIpzFzCxwDuBD1vnu6jaWEwt0hwsGxyTocGAgaDebV0Pl+
aIbhk2AruhRVLHjp+uJTuUQwue60h2XdLi37hAXS5NQzlfRkH9BKrfwzPXghG7VE9Sk/L3Map7JU
0XYmGgha3Dfnphb6XWaps+T4KLJI/jGlXsf4eMi71AKjisfMzD2CgtNbZsLdHKjov9+al60zunpV
L871zhwBryPwlp46KnKgA+6n+GHBqSaEZ7qWnTiouDBo0QwbyQV3kqSdXmV+l8B6Uv3ZvABe2xdo
EHlEJWGWzSfilECHDE0cjpXisqnxJjhh0H87QDOt4tCX2WhbmhuyfSKtVvl3pKvw56b5HL0/OGCR
XLJMTell4AqDWiibNWiOh2PaaRA75mmesbDad7xxKT85beWd71175d+TNSXJzzXP4zYzinQxyDJX
HppNgH+ymX3qXFpbcn/4OAof7H90/JLl8SGvMxx6XtRt+f/GYsE/AhIvwxWl3LiRv8Rb9vNT5VHg
t+g7Scak/mbAhgwLcXwdUsFDCJlajgBwLUiANoAlkqAPoUyxUX32IADxYySQ1XwQQ6OdQDJEyqLi
zeROipPZIY7hrWYSwMpK537w5ibD/340TewH89p23AT1qgIwbdI9bIoMa64x5mXtaWYItpM9Orgv
pFX6Agsfynf4NpABQgHo7xFEGXZKoWD7tU+6w05wpUUpxWuUvdHDomJWymHIx7UglMxZ/uyzEETO
fuxVMuSRpPPKHp7VmluIFGrM+uFk3eAznrkJrX81kCyjZ2A3XdPQYPx9zLcp3hW8EMZBv/rG/Kem
ElGenN4yxhAr5CZKKLtTkIFJRqR/3PlA/CEnAy0k4gyJWLGsSsSJ7Z/hI2WNoPYa+OGhlpfGlxMO
jiSPXRb9qqzgsS4aMoHYGmMZYqMSX/LWKGljxg9pPHBhZomcvZYHNHqDSyVY1XkbUNwH4j9xwlSn
zk5PbArWeYGojWgJZoDnzv/F+keBTxn02PHUE0bzssAc1J3SaBB2exa/rZRheGD5HuwnKEmvUaXg
J/n5p/LQuJmAYVytCT45BQK52F9LB9Qq4YtAIknZhKf9FTgGyvsuuBpPckfNVwU5YDn4hc8NIBt8
QIr3ahGDw3MNsrQPIdl3j+H6rKJ/AKyLIq5HfCvPVIBX2jr+ekkJPoROAycthLxiK0lQVGrBW9yu
gX+bTN1f79aH5LTXnEGDr71wXlZ/Lap7knRKnNIEdpGK34q6krSEF3wFvSylalp9haDhibIGIQeb
ae/uY2flerxyb5b0hyXBavEymX1zVjdGwGKqMcr4IQ1SxtQvd4m/FMEU0N9Wtf1Qat5kX65i+IlS
qarUu1NKDnZtlnAJjS6KE4vUhxngEJhvDsHQ1OZyoCn/iJheEAWrBieh8Ypv3sCvRlEBUXO5UuZl
c4VUqXl8fVy8WuGP6ERpymOBSSozK+1kCUGsExt5cHcoKYNUfIK9Mqok9D/Y41uxU/eLlxchrZfa
uVKiWd2kRl99Ec9CCdnzjCwSHK4wl/ewCGlrbEGQbngSv2O/BVpveRBskxKa0eARi3EU+s3WyNrZ
Guyzxfm89nML6JmO1Jb1RnWMYXYzEqGJe1VVL4PxRI3t55NZ0XCPzDIKnhE9JRzPFSlzhNUBtsqB
DwePI8SKzedJaDPYs4I9DVSiScbxP9NtOUqFDoAwLMSkmjZrpwdy2PIJWplpaPCGCYiGK/i5uqxa
oin8tSPSFJxg4aIA5kxtdrG31Tx9GiXNtBxF3c6ioRIgTEG3XbN4YdB19YfKd+1XLSp7OD75kBHK
EtnpURimyg5k53Gj8qhy7lUtNemBJernrLZl34RiVWlWGU7bY0w1R84j8NqyQJiSczImipnoMmhm
ii0X3OQIA63HK5JiHsgXfEQ1jZg2RSKpTfOMXD56KL6eza4aqNPh6t+ed9rXC8OjQ1wDukW0QjEW
SDy1E4wYmHl5aByASdbtZ650Rf9sQN9GjgLUhchuVQl8izT4L3fT/gKPVyi6RVkprYapABug+uMw
WZh3Sru/DKn9Rened5Tst1967TR11USyo1XklGyePbHH1ZhPDLZYTfzgvQfKJtHRl3UMUPWA6tgi
WTSfOyx/+fvqQdCx+LI8VsUiEx+Bu66GjW3/IC3oQuXLoLo1kw+7WT5+zHw2zPFyWWu7o4c/uiQe
PnpxqiFc6VpGLHl+9YGW8eanPQUyYmMshLpFiFpdf0YLUWlVjcgRVeFfJEwhdc0Exvyj4FzxRoie
1Ol7DkcHSM6PmyLE2/hBlvAk+IbJFXPi7oBeTqiMczxrjkJbdRM+5bQf6zsfCOxyJ30y/xF8hwNk
whjd5d5yM9rO6DoV2h5Igq/cpFjugApqMSf9TOXbvB6+57pGEpsGjQm64xkIftMdn1kNz97v/Ghy
lL7HNCIi+V13mgtR3FEHpHxG52no5GMY0E4IYotyRMANlUNiQv/9FbahV6IF4zGysK1G8b2Uqr9p
P/cXuEmzgA1azSgffcm459DmL+APeaC/ojZba5gDdaxHKZu1bRTip82UBWML8Kra/Sd5ENAvt6bM
4+ocylLvPmOdYuQF9JYVwlnSF+ljOHrovsM8wloVO1SXbYN5RVcZisztbXlWQIfdXnq/UfhvO5br
Xh5gGgK8TrtQHRUk8hdEEDi5vZcC5K+upKqxBdHR/e19PKme3jq3RjB9F9j1lJz6f2tBqCosjM86
Ar17/ea7VvGjY5LsQZydHAxNEf3PASEeq0vcRG2/hWKATJEHU/TbQYosTBPu3vKH9Bv5yBr4eac6
bmmf3Jgzj3498M5Rh3/HbP1ZSZxc/SRzy//tpRjh8UsEsND6hRjFzMlBQpOmhH/mzQXqRUUbnSij
lZJBvNSE09YUhBJ8jkV5atXjOaTOrGUrOCteGGthHdXM28K6usLGNNwASJStTR4seds7sK955U0N
lnvb0vVuP+B+7CiukdtR47QoElCxvwMtcya6bTDPPaB0rPwH829FgGm5NaUqKAvBsEwtdoiUFAOC
h2oMfkrMeu0b2GrwXt2/XTpfxrT47qc22MlE4BKURrk1mvBAPoj5iFudw+QycmYXNeZszOH6Ng/C
td8rTT1+Fr+L1zR8qBufkrKUXHbFmJ+qQKTsFwhHr5ZSYjVemy+KYUjXgFHBJlhtqJXSr9iRLfa6
toM4+Zela4iIYhEsjHNlGzWRiRsJUx3B4S8QVnvigh4b16nKKo2AWXEmLUTW7rbYrhBAN7rr+LfO
6PGnWhQ6zygWFXSUEcwxomXedY4FK7g3BUcagG+mVtLXoVyoywzMtda1aknrRtgH6V0h55YLzyFE
SyNgMkHXVCTeo4CLncaMcehKAxoCMDx4yczoWg8QlHgAezpcMLHnYz2KtMCyUljbi85kpmufQXIM
YgGONLnlNa1RhBOEJbuIGDKQZ4baCsG8vjLE9s2Si99HPuiUWfJbmzjtykJt62IaVOEWMCi4fQQA
UBwPW6QstCIlVBYmF6nvgul1/u08Iwfq7ckQdv3lk8QAEykMWAarKuQ9MqwCJK30ARqAz80Jkg7U
hJ91YVy9AWVlx427WRzCQdSbfQv459/IMQEkUdCb9MgAfbv1WsS5y/PxdTwYOaG9YFLXIH+ddFtt
OqZrvVf10WHPHFKGNgHSXqgh0LYLSevOVXeWF7mmTGEvLX4sIvd0fEhg3HytAggFjiTVtsLz68EP
XIuO9U5zNpZIS26x9yLkspeg9i6Y61XJu+yKucPrZFhkbjV1cUzeeJdiE3mG0STDJKlb9mAGqJ6k
mQs7+1gbHVpg2tn9NTQQdo/17CDchIKfbHVkmtR0wJ1zFnA1zmm0cAaY+TYu5MDYaLCU+Gnd5K2J
G/C12bGg14blr688zKRr84zrsJIKNkjBH6aGLFmcuB9wvCC4prdoTWP8duVTVChhNqgjh1rX6Zi7
9np2nyS2u00nZYF2O8cYgtaMcXRd9MB0SFzle1uEwTzM3mh7yF2eEi73jo3i3rBWSV/gXUa+sbdr
+D/7fWTIzwBP0LPXMsm5rAfUmNBA4xnOLZRxpp24qCeJNsSiHwkRxvuxpD8IKYV31aspt9lsuZEe
gJr9dZ2EOwSNFUfnKUIg44Lm6IhzPBdbygRblWBEJcg/KINv/K34xIak65YwzZU4Xzlc2Io1/Bv0
dPreGLxTBxs42dpcm2LGio2ZjwQYZ7b7IIAbnS4lVlkuGR2YyWXv14WroWHzR4/Vn0sphiooH/hS
b+t47G4d86nyKvsra9omB4lgcoavFxYJJaryguec/yKMZ/qgpFevIuDFTYLCTn4F6jhbZP3Ql1NS
SZjoSwQYIG/IR8n/dUDcj0wj0cPtBTsPNZwLkyFh3aPnPY5fsC4kZrveSOpt3CsZkLGO+QavPPj8
YxfSecIUEIFSJDdHO51f1eAV21DLpw5YYxXwtkkIYr+tLV5nTCX5Q0uX3od90s5F5Lwn2TrPTg3n
pmlex+5j7TVuWI3lNAUlnNfaLpD5DuoUEaKJPki/R2zkENJ2bfUaDv08H4FK1ZwAs+MGm8BTLKJH
8rca6BP4PqGcmsm7Ba4+gr6KgZE+6fujdHi6j2a/AzmijKxb0fZykxW3hEIG25VvTfadDVG0fHWo
5VMWyxKD09N/HRFS3Sm1rfbYdj0h2I1ZqO1n+o//cJJqmtBGoJn27WoliF4U4fzKqcNG4zZqKRkV
pAsnmNhas15re4cSytY1O7GSSsRsEAQEZbMdTdN5L/MhtadIpZC6s1OXIw5vH4yOlRYGf2YXMDBj
8QIEdVqzz2FJsUVtLgWak+Cdg/WXvWDhL7+FO+SyVmMDVz381zAUdvzoMz9b5pXVfX9cI4bGqTzT
4NRVeUjyOO+DgCiPrW1bVdR/fBSmuSVGhIQupBY2UcRSyt3JCNC3Z247rcsWnUJnxMOKLDHpgLi9
ywykhq6zFmu8JAyJSqcJ/d5CkyTzorl41rB0xNNZjFwF436D/PY4YhK/Ajyq++XXx0fhG/+p0qWC
csT5h3+RhOciNt6F6zpVgV2U4WMcwCuFlXZUgtG2lC4cfe6vCEsxSnPRsAhx69uytZqV6WHlBFM6
1Zx3Bxrm/JXG0oN4hRBc5hgtvdqxZ+W9+ot8EZHV2IVHCz8Ef8ORyHGzH034xFLZK930YonAtNMM
F9fBhbuHND/pAX6yjkEBC/kyh9lePmAmIZjp+oGPwDLgXVj1W0BxfuW7zLNfct2DZ2ZGGQ5rH25l
5cCPgyhf/UiZrbfDxM9dP3/nF872fYjLibHj7xG0HAaKzRx55a6zOaQ5iZxSBb4Ni3/OYIOkD9pu
S5q6uQbpJ0Mf7CDgZOm7ZwdTUou0QUIX1IkHhrdlcgtxM/HRgRO14w1XvwhhSfzDT77y4fIKUhvC
vOpCDWXThFtepSNNtqX6HCp4I6iLChjHREsmqqt+4edHUXqSiWFrfz/x20NyjfKCe5c1Va/Wee9r
+pVUyEVN1lfdlPET/2OAfnO05Hn/zfyMGCEKyJXi7pbSHUxLEY2i1sEHbnoYgTCFH6wiNtV2/Who
87PuO2+dZO/ROY/caJfwIdK6mFEeftKjx7xLbNvY237+Pg+oKGwIiGperC0SKZhyxmhUIwz6VhiA
H2slIeiQZDmkMXxQ2aepwyAnQzWLqZ3ZhMvvO7US1P+dwAyeonxlsmOQan/EFzCd+VOLPj3LrSgQ
rusvBUTOdJ5wL5gmEyw/79as7tJ1d9Zot044oU0/Mjhoyca/2OKqLmHP4RdptJCJk/vx+c6DWJII
+KOsAndLmKSdDfoTyXLWM4pBBIWMKNANd2qOiX4QiNPjrG3/0yRbtE+zuhIMaqQ1IxGbVmcDmCzE
jNaI12OpoAtwHUVAvHU4rUaDLIEN0gASvxL3/na8IBu+HPsQeffsa9tygGfIscAk2jb7Pk2UX86l
TqWUTKbQsIICAQLhr83o9/zTD9aGPXICY8iN93ar6DZpj7KMQmpNtrdlv2AyojOtKw25gTB9hcVV
dITgHVAy/TV3OFvYmvl0vIxPELOf7GGzNulrgQvbmEPlegYF7Sr73QqMIEx3Oz6OREM+1RQoNJwK
C10Ozrd8GPWtyVL1chkyfm+MtcFVWJREME3vA/5CC77DtqVe0jz6q/0PdC4IjSq/6XZVjMVCoe5u
luEb98n81efiItr9mRs289P05UKMLyIESB3HvIcNVIQpcK76aaOaptJR7EmERVuOZUSoVFPUUzKw
dPsgwVCtPOM14E4A4yYWvSDpVVbKneMpnALC3mwxAvTDKWzOnpxpFGTb/r+hoxBJ5O9fprTIKRKo
YwLiaesvQ/cGgBuRyF+RyhBQXdv+hoi92zPXCCYTjvP6cn3h2yd7fpsgwPEe/ja4clV7H8cuDScU
d1pkbxO5aIHTcJNk8J4qIxv+Fb3yzOfBqeva8EVtUNWSTJ/FlDWC8OuRN7+eylyar2sFxeSD3n5R
E7KE89BRR4XWRXwn1XGyWHsNKW/cA1Rc/4EWhboKl7dCL/qoS6CCOkH15sfwrqBzyBAum+U9VTyi
0MZgI4mV9Jd7PKhGdL66KNcIqlrqnMvib8CrQtTpm2G2i+mn1As+Wy7QpGRRQswzFFpdtv0SuEA0
tigmK/SPYFw9DIulJexkEEKAZSuGj/Cre/Ub/JfLsXsrgHX5HYLRYq9veecTmfPsquAoIkewrmNs
HgKHCNCC3baQECI4415bR0oYgGX86B0wiwmoE8VqzZ3HjEwCuCjspo5mxE1WchyMNXASyqS5sn6i
KiSfp3ORmpoeXFGtnrfNvgdhhuZfTi+nBPl+9HyBefQrhUi7WXYeHT7/0q1kE+KHCTGRkX9R7+67
BR/31lt70HoDLh78io2UsAv39C6JEscORLcQ/qDxIFtp4QJdeSv+ADKpOMmS5fje6lCGNXk9Cbhx
PwHs76skcd4/KmVM9MTuLrtBHAGRzFzqctQVnQlG9gxT1Opx+hazTngws6wus854kgKEUd642SqQ
UKbUYnfkWyM+PsXNXprfuV/jPikd209rKUY5maIJJg+/mSsuUO28pZTGcC/WEPHu/kHGgYe3HpRa
Mqfz9H8mHpTh/78OJKZE/wapUNdQ+QQSAk0g0VGw42hgZkOJ2/kJ64O7zJM3hgl1w5mOiOxcmDn/
E8UFbset+pkXDphZqKBN7qIPubMcD45Sg46wVz7LZW7BgZKF7uFiddrvjNA4FaLqK+8OpF3GFUEy
HM8OlcmjzhfF0j3YgTySgNvP2U8rilnKsd+3IuXGJuX595FATA5wuMfT0ofdrD9fon2Af0YYQvWi
iFB7aLBcK22G7TS7FrKZJY2IKKYEEXuI0mvozflEIWFlKt9lBB7EjDvRczYEin1OOVyv4bT6FjtT
Aiok1Rs4llxByG5FZyC9YcX0uuIwZARgdWQR2mw1PkJojvhJROe3tS9S7RRwQqRygo07BzyB+1sr
xy88zmCKIRCKEHXhzihgWxVome8MzCxK6XmaY2dfNL11+U+hiVqayrQI0t8WlbRLO3/VLOPoGstH
z9N3mIhZuVuGkNwryZw+BB+zE2tKb+gX7nSqOMN/zg8IU5sOMKgu8iR3TJXxOtZPZTVC3odAVPlp
NCBtO+IOnbKdbaLWn92678A7ASwdjAgAq1hAKFG1WLW2aD5x0Hh8ZBZbYhPDWgWG4SaG9NdLu3bh
xVK/Deg/u/8Vvx3U8MfrBSSy/5ZR9H6q3e2+rdgOrq2jpuEvOiq0Glbp5A2h7qJl/Xtq6mBr6yoz
rO/caMglbXaIbPaU+8BU8V0+MKOUQXKOv8WIOZVd8GzqH4Z3pNW9ZJSnoWVjllES2WZcpc0lo3pD
57neOPgAyzUzDmdyDR6GE7U+yhYlpSuQxNz36p9+MNb5VNQ/rbC6HvCjwW0WMMAWna+pbCibWYC2
/KPAgeG9ye3Q8nwHdWtHkBMEarDsCkLjbLHqejw1yLzACmdp2SOPVjVmMhDXQiTv1uA90Oyu3smc
aCmHW/PdyxGUJqorUczo7bNLKUGn/FJaUdq9LS0FUf8ffirc8YgKqbFoBMhxtcgXb9YRfAyHiQx8
wk+FxOohEPmycQepO4i4ATFeBf+JOY/+zVys5WBWLXeEZAiEMi2w7xM8S/XcANP7rWQdfshH2pD4
rt9/k5lXnqWYgNFjbikYKmjHVxueyQSOe7809tnxkik1k3qDWA4+eX6W9dNF95Rw1wL/vklO5AuW
MZYI9yIOvMuaXfDurn56lvDuTsUimLdVrmOS+nV88K5DakWYaE3V1D9YiZnf+EDrUpWCSXc30HJw
Cx68kkRFaFHA5WjuvSSMeXlMgKJQKZQnsKh+IQZ6mScii8XXH3Rjpn3M7wjz7XGs1edQ1uayYilW
T7jXv6QWLgZga0637xSpvyimWxYaWsx+cFf0pTOsFcFOUEiRA0qfjD0nwyLfZzvffABfkabNoPxq
rquqtT9IPCc3b3oiSBYGUx+1qQEcP1l/VCGociKia7UYuYwccnwDDxHYWtRRdgUfK+KYYV1bPZTn
DAEJeF0WjEpQ4LeaLnihJsQq2Uuui0cbpNfek6gYEE2lqav9QGlgiJuWypUhfAX+jY0M8wvwidm9
ZiiyU2Hsa4dFtctO0Qqx6uVJsWNWv3LYn4M2WGIM48IRORlEz38TEc6Jq5L2VUatJwTVxBIdAEbq
2n3lTfEA8lEqJZh6+Kmm3ol/FN2J7tEr/VunpXx8mLYT2NXrHrDjgH/JKJZYpyotSosPLt2Gu6wF
5RwD0y5y3QQzs3xM/V8ubG+8dkA/InpDBiz3f5jwa+6dnWRbZ37Xd5u/SU251mjUqJ/s74u9uLWM
SMC3gExgqE2a7szvYcPwpJlEMe6kSE9QKZ88i41HcTwv+WFcXN4nL8PYYmhAbgiiKw3qVA/ahSka
bGWc7DmIDtP1SzzJ+82lwjKPQrKHLU+/GeXb7yvVnMtnJkPbsFcvtaJ92Gq6qXLzxcv07XNAbeWL
uCVe0JhTXNVlQAY9JBlfGLs8ZwqBSGqZlnZ7JMDBvFgf4g5PdHzPalrEBiInRhkdCWsGWiguI1Hz
2anoMPzPzbSnYG68OztPO0IrObdNaDsjs/gvmhy8h1dfFqLX3sTRhcWmnB4mO/pVVRuQtdD+NQdI
bAAzl6KluZj57WBgc4H7ft+ZA9z9dmEWqinwVhzuYHls8uC48w8AwE7WAsO8ACtec1WRMKWKTBEV
gnU1hNOgjHdSWdmFThdK7KskuInE4v2hjru+yg/l3wjgW/IvAfHUBltdAV483tVr5Jv0oG1kahmY
xTJhJqRuYmQ18jnNYuGlRT+OCUeoBrIeYZyeXzTihqb0CFM5jA6zTlsSZHyEXfwS2I1yeXepjjpW
qFowSH1cKrNCdY+wMWHfpuDDqFmoKjOMzvYt4RPPbc1mUNkqp6WooGYr/qMTvUGQ94HJm+bTZJyL
GNEC54DAgwBZ6xXCRN1cXO0/0aH++9k2T6WSkfGIQARJj5mxOQhAahrRQFysoCH+hQXlQQZ3ey39
R7VpZIyMmpsABPm01L2MzY5uaK0goqwDqw3QuA+Td3nxgSTyHeGfIVK5rtv6o2q4CEZSFiArcwVw
HZVpkxb3jqOc3+29pWahcc9GmIA4l92pnebNSS2Xr8BvZph6WatyS84kwTg0yQdem2/sit8767+8
EGBL3qODjOaHKsDvg6xw8jGpCXBB9bGidLVYrJgj1tFBFra4dXiI3sc0jN0ylOSz+6W4amIzKD3I
u+C/2ddYj5XsAkqkwb8geqGMh+eCVr7HyO2ufHfwgjjNCh/dcGIpp89+73ET8NiEkl5I+qR4lSiX
mwqWlpkSXak/iG7YXiJMWLp5d7pOWU9nbLemlBXWWEkDefSAABKQRgUuerlPel+Tz35v7p0i9FDQ
zLC7ohQ78SI9ELcn4/QKr54IJLEhnStzHtg11glMH4Uqjppmtdb0FOD1KK1YNTVxk5cTC3W5oedw
xin1M7k3NRGcFcPhWRxjGk9o3S2xzAO4IIGdDUxVrdPMPG3QUdGUsoiFePJAqxzbdUaMprnRX7gC
H7ypNphSE45jbBGO4O4S/bZPshGpaL8+XKwKvpO03rK0qkcEgORB87js3PiC1ydqkCcXGwtIqHDb
uW/jZxtfFffEm9cEURO5zWo+auLo9yGgVoHG4ZXW5s3yAChu0+uoeH/njM/bpR4lZZGdc0LFB2uo
8tjWYUWFhXtZtdmb1Raic3naeeKxzyMcA4mRpN2pMtz6dY+DrHaOaPavqiCqRxs6zEcptbSwa32+
GRrNY+NzXzea/Rmk8dXFi0AhWf6wAoS1BrDhbNGiKCjZClYyukWKzPs8F8g+rRoHUwqBXOgJ/Wjs
ABc1AFhrbxWAeHz7NQC+PlZkJn1jsquXrcEEizHiRMrSnL+eU6jn2zs8pyXklqAPyM3d4sbX8tN3
lg3zpmDjNLtdQIGmWO8z4g9WnWOnFMqoWEPZ9wD/OadoAieZz+wmE7SG6l5sTRyJr0GuokjZkCm3
9KxPP1CApn/yidzZv8I5eiCvnE+94TlAeCwi1VLJ5lxGuwTmcKakzgRh/3p4mGvae1Vdy8ryFgQQ
4milrBx+IaOQJ6flZa8fVNmn07DnzbAoU7i81GfszgAqKZWGecrobg+2qTbXVtCbW+vG0fzcR5Df
5cHsTAlYlQ73e0vGzLUhX+mNzS4ABzTIg3UIlLDxBDzWUtTrVqLJVuVVGL3AYMk0w4mOtnh5yI1v
N5F+pUeAEKtUagLpyn/YfiOkBjoX4sXNa0S595IbpsYo/nb5i0bsFUrl9eHlryPov79YQcHCqQPA
d2tSrwjDhuhEY24ESCAav+kompihurLvSTEwx16V0yHvKc/FYv9GFdaQTkEFdKtEY443lLAxGuU8
HwKoItJdWx4X08u/Q4h+mXg6yOvvFx+pKINstoNYEovHac6bxeYcMMqUKfqrji+R/P4vTUrYDsM1
Z0kyXjnNY5MJW4PGAxW5x5s9X1cA/DeaCgu2DhAag+YjfzMbOOOpEgZBiQc1XqAS9skQSAdUXOuu
U3aSEbBgmQqR3swk3MDcAwN68KxnJafB3S/qG41Wuf4hdezJ+jkNJfx2ROgSIllWsx5Z5WK/ASBJ
ng8Atk8IRLxmrRVmScUZGQpXcA9RR1BF4FB8xP0zHBEnj+pkQqc/1PB0elYtr57cyizkiJje9wzD
FVeJUWcFQ4fFxvGds5MWn1QzlKFZ7Nm2+L0qjjy49ZN5TRukf2k/EQtm4TD23zc4XnNBzOfz0rob
1/TZwuinauPn/FXt7v/pAyiqCvUcvMCz3KjbE/gTY7mXWRGWy9rKmLwDqt8nsydLiR7VxCcJ7Q1z
b6jDRXh+QKZDFaM9ufwl9k3pvS8SytHH+wQ29mdn/NNkF8sRLy5t8h7QLtxSho9EIiw+hw93gyMH
WviZpDJP3/Qz283m1X1hraiVwx9ms2elrqXOXYdOyXEHZF7p4y636nQFfGTbpkM5ZKSrvu6t540I
lfd7b6ju81iqvJPiKI3YPaI75V5DpTwHDgtjH/LbIySCVHEr+H21BadwZ+ToljxjkMOiv0QcJYEi
4JjF3OQukqtQfbdOKWBN6LpIF4SMFr1P+7lN60OwlXZKq1zLg4TRWEvPwjLbVQJgucYOe6E18uhA
IxEb3VO7u2vt/DmRjp2jbTAV+rtm6tpU4AqBhf5Kb1cv3PjS1fHVhFbC4GMQdbYiVDJf9DeYkrXb
555e3G28hcOOSD78QQwptudPuCqJ1qLtMKJFBIyrQr+5TxdpuzpwC6fYkybjHfh+ij2ShHw2Tf2N
l//tb7qV6l1dglo1fJQSlYXe1Tjdt0xjAVuJFhy/z4/VfWQ4zf3n5iY8OR3Pr5dmjZAWhY8jYmZS
S8UIiN4IWWjSWsFMqMw6k7TI0n5jXP6/0zfMXmldoHN3HsNdmElnBEZIQCWg47AFYZZ043XFHZsj
7Lh3jsK4r9NPtn7UXIW0BWOntADjBJ3rNShbx8H1a0JGTLT6YmEeR6fAQF7VZ+xdkdQj/5aFlaFz
FlLSuUrvQhTJFxRhtSQ8dT+Ur6MmQh9K2jmNt3ukrGjfSavS0d4Vfs/bC1GJSk/hgiFw4DwoFgUU
R7URExKwR1RozyJ+G1oyu+jpbA35Zk2dvpAY5qFrb9laFVwgRtSr0M8cQBr/uxD9VQPhpM4p8Wxo
WDGby3LRGBNm5EdGqzsTcm9IrJb03z/w3JJPcmqq1+khJVV8Iep+e8wgnxC2r8B8hpIAYBVChwwA
xBKZXJ28iH8mBUfP75SUdxUaCd3/ZSV9pP13rzEJ6GKCPAz9yWKS2kyxc0mO+XzN63edgHFkzc8R
S9hF92eGgY29/MHtx2fOlotJVzhmZKEaaK1KJvMWcI4GwpbICFAykEl9010VbroOv5u0yv2F6S4A
1FmXIy6oOcChODrX0Btniu9mUZcwSOPCcG6BBlnmDPZVqrXtrW1CIAiMGEfbyl0Tavrm3Kdn1aBH
S6OjDSKDgrh5OZ1D9M60+/cYsWQ0wdn1t1OM/wW1dJyJVu/wSsusi4dW5uNE1HcRRBqlv5fKygtp
H9yYgbZHQ68IPd/jZA7nv8MxBIBK9ijlIAq/6xrsj9xva8s8rrYW45VEPKNsLFM/Rt9GWOafkcpw
kNEY5hPyh/dps+y4ahS6H8+CUMCO4w9qWtBpWpr8Umz6ie3QZNa3nXzzimBUyvpLTpaWdOglqZAk
aCi+PRIdPkSbSpPF4qcIFfIotaZ9sikDtPb904+AWXSDBjiz0JXY1SCf24UCBkoLdiNmPxXdbLL1
p+XDlVnGwlP7L9pqEvBJZvfQBikErXRuZBl9y+SPA0NlDJBO5A3daS8qRWJx2VvcptoQLZrP90AX
1DMDH1LOL+BP3zyXjHrAH9SK4iHWBpEE7ae/1JqjqHhGudpz428GIcNHq7vCTL9DUw1Hy6r134BB
tBvLL6qavuy49f/vTrZ/DlN1nskqC8wFOQFmOfbdo9DeRi7YlCjU4NTcNHull56AC7LfHpj0NMq7
U89oK8ZsSRAn+m2ZEYFQIv/nn4bg0/1WF+SrzQpCRs+9Ecx67GpxFfmU74CIRtv6yITY1UdDYMbF
bU6LOc/NxPMR7J9/Bsd9+26MbagZcXyl6ReUaxviPITgXaS2rJYXEOO5MBJKkUpXrgsNTpnNqi/n
Kz+tNEtkYrlIJB1MDmJ9OEGT9J2xWJxZffMXsH/9bXmBBYEatrK1N2x/ZD2ZmcVDgXhh2VleY8dQ
SEQ+esXINlqFI7IRRwt5RTrunZ0Si5HeCf0VlkvarURZYPAJ+1e/Q6nYvlYT9NP+meM11fdRuhnP
zP8+VvGh/18yoRB6yrOl6XK3kDZgqs1yY+ps5ZB8PL2/xwuXFQLS4pT/N+BVCIlLBoiyNp0gWQfl
li/9yZPH4ccXXZC5+3lXslRIUuWJI5AkqAYNMWcZANUwrfn3hvSMdFBmLZtJHr3pEi03MNkTMIP0
WndXNDEpNYwI0dQ3I9pxXx6RP2e/YjOv4PyO+hLGtMs/05Q93zw99u4NDR/4L8guq1QfzRcW4xuW
x0m4K44LRvGTH1ZhWgmSmc+gUnPl0rZDnGGF0OlSG+jseuc/3zGYckk4gXgDH29VkN3MEU0mSNB1
PRYcTsWf/el4B9hVHQACJbQ5mnOd0vKsdyhO2p3fI/MgdsCYY1rfKPDZgirkJsxg10xoFvgR7+ZT
4eQjrKRJ/KhovNUX6P3utfinhxupvkFkojzlym6J8FYBqLA94RSXSKARne2nnGvjvZrK7ExA75D9
n5rDaQRfKvhB+/IUkBfINnri8xlMbAbHzA80Hwrj7a16rMOEpIfoiz0/hxrtDhk8vn7dD+h89ci/
fGjSR/zdz/TFVnuZ6dWXujgQTsGGB18VhDohQ9iGtq2vl3BgEm3pRDJJ/yNIao48Svi7imR+kr8M
DpP6hNR2Mj6FVfswYKQvhsuBNKkzAv0kSHoy2s8Eeox5ZjHNWwjvdPlPX6fbWF/IoXd5Lfll0LeM
D0OnzsfTH+e5f9FabJHVmyR4ywatFhkHxWRCZvPwHmJi2RwbKs5MrZ5XZWvnzFjWWAJnsm47asOG
v4mlZNBVww7ZUZoypFyMZFDAaGwFzCpZ05xKx4P7OHdjRp778pG7Sr/CNPtN3O/CZZwkTNR9X/3z
Fo4/p5zovVFpqUgTYamPidzlPBe/IOSq+kt9cs21hNhpzSzI6etb1bb+v0Msu4Tbj/vEFM9zJlgk
Rro6h5ZXFkRmD+BipT+FbLl4tEUEjzAhdGiukdk9gDJHZ/IEX/IUjERFO4T2NFd+dmCZOSIEcgIq
fDDwMwftquwNgpewjz6/VZ1yc10k1IWe8pI6dZuD6puFMZA/k+gUb/wjnvrdrkhxkn90komV/pKo
tqujksqbyf4HJbN5b+elkfRgrTgONStghNEbGhdIHwM/bq50sFN0EfA2xMvg8E3guQD6VfUTShVJ
rY23syAdH25S839tmLA5mW/GCWKsJHHzsBDmtfHbPucsEuw5j1AAA6awY5FI3qTAuAU1qMe916Ae
eMORiwKewlhxXHLj4DVUU66+yKbtP4iFvnuU1trTGYjNbl+vgoZ4Fu5x9kNSBNpjdSSr/ydo+IWO
2ALL4gR3XQlvDt5NHjNfRylfeJsoSWnF0HTWCBjg97RLJQJ8XVHfLhmTrHM99vG31M0HrcpxAZMk
l86/cuK2V5uz6L168e5MkDIQhzEANUH+p2nRXTY4cERASjmWuX77iL2IagSe03c4ScEqKtLXdsH0
4w3zxEcPuf+dsp+n/nIN2kYL5fANsheaM/5rVAPQcMqZjq7Sm4tMtLCIkHGSqOCgDvJD9WclCSzl
W71KxbkCXs7rLBErEDq9PJDncpYwGF+fkfDNOkdY7a2C5t7M+Q8ow7oB4hqg6/n/07fko4qD84C5
SrL4C+S82Xr5fK1i+XIXEd2QciPUItmGOwRoxuUs6bW2wMTMoVjpH5EgoSaPHCU9YGhvPz4O2uAB
hJAtqf5dPBYFjPkxKZ0+xY+oozu5eTkSuvHbsBN1eGhGzpcCx0FQHByk3DHZ0zr4bZIuyMDxrTZM
zp7WgsCgaWpyl9xNRhW+9S8qbABYx+O7+lGwMlVdljb4otj8GksiM+cRzqtv3U0ZDV7+pfyh0HUU
CHv1PC9Ltd0DQMy3WXD3nlJN7+06K5dlfp28Maln+WhN/QB//bDRVZsEXBZmZ9K6thabQrbm2h77
PQqL8s8hvw5O/cA01JivwVZ8IlelzxTEWsRWtKtjiSHibJWbnDR11htLxO13lV4BCHmE1Kkq2Kow
gQ88O0s+H1CDoneJacExurluqtBqWhfEAQE/kZq7zv+oZeJFusvUYkGZWBZMO0qelMJWJdGSKxSq
CRZaKNzUtAz+F3C/fJEPzvV6T8PaHxpE+F3K2hHSF4bkqIlO5CFyELiTyMysCrDhIOApDtrDLVSU
OpMKAcKMfEniEjE/PQ8u2QnIwQl5tRkHisqx5+YU1BTyN3wkkJ+zW69IRor+dCxc28a1QW9uRZ7p
cv7fSjH+YuWDD2/mA0zq02FmjOId5OMI312JUMXAMrZnvyydgBg7gc67NclVJvKJ8OGQAmbu190k
0FOduFRYM3LmUg0/TMtlRq0nrejpoygy58x7CUkddv1KAbj73UTCrMOXgN75fpVeK0sXkHZJK+I/
McuPUz+3CxsQiRf3ll5uOwv0388cRgqENFvUe8/Vk5HL3QjPEM84DSI6OoBtrAgB6tGLX+LbGfzW
EjkEZtU6Su89cgn3OCpwV0Mv18yWN1CLa4dYZHh+p+zv7KwSrJsGnFqAGviCjmc0eXdFBTRyviYt
m4Ig5EHRa5B4FjW6QXnuzM46ilUeGJ2FL8tO6C34T1oQMdpHDpFfQ5F3E9rRSoMWNaNCfWL87O2d
9Mz+pqdj01WRbPQAPr1Pol1GrF8J+BEYyztpfzuNtUZ5J/4d6Cw4TcvWkRnBcRhtUGCuH7Nf471Q
IWNdYTLa4ih6FKOnrCsfQl5vjeNuR6Xt8e6m+S4R0cZGRzd/vDAnYepbkhW7bu4CnGRdE/BOYrSt
oIYWZP2KqAsLAoOz6wDakrY6VchrUZ/3Sjl0/nutyiTWzE3dW17Y7KJWBzSIHJTcc2N6aC4Szqup
zUlMTSRmCUNCOyq0bBYMYiKPLikkt9ZqNrjvufYmR/hArG46IfmGfVyYwRCvTzHDvo3RG8vCHd1d
WkAUYqAavPC6jphj303f/yQSjvQKvSvXbvUDgsdEDggSvqgAmnm7Z6bVVh7yoPdPf53vjPRUi/71
SIq4wPyEKZ7DYWYwPVisGz/dwY6sEfZOgrAJEJsdfZ2zP+dBecTSjVqkk98VHOI2Ho2k+0AJEy4Q
KKa2FiiRhLASmP9yOOIt7aJyHxi6o6ver+tCuz5pa2dzwmcbiMnSTm1bWzRB3yCQukSQC/1jzjv0
f+8QktZAKpBT3AkBx5lxXUrZGRtlKvk92aXCjX3enT+Fvgy+DzQ1c7J4jbuos60p39ZaPxmX7+q2
xs447m4kR4DXK9V2rCPm4tWCNmz1Z9VsezGIzqAYIZe13HhC7ZDVhKlPPad5gzvREP7Wdt55BnGz
LpZZaIHGbChIM9QUgNlDLFGjcsGfaO+f/Twf1WzEQ9ctZ/7xxPrP3bEo4gL5eFXHczIAq7CspMfr
Jri2RHPwRkv5YdwZ3pZR1HZBVSswazz98Ok329rsj09xSGDCw8RFdsgEIuT/9I7vL3FXE8wUaS10
Z1dTFcxyEp5ODTxSgUE6A1rxlKbN6nwdekt6hVOSAbjNn7NK0CQ71aSss/vnJRjxHnPUu6t8aQyi
phEmcLYQkCw9FhdTBD0FOcwPkKJt2C0CcNipPR9iEA2GXKqMDk7uUGt6ZTWNAW/mQ6dY74DEzcUK
DeOiqJ9tGZT7iioZF04rjGJVHmhWVPyQhkDdD0kJF/VPCd+8qLbj1lx3gAdYpNuYrQ8/pzvgQlMm
pJDh5yKZDdBs0Ppvjiy1cVATk4ObcbpyZr70IFM4ZV/KukT8BuyNrik33S48+r86KVTKo4yVKRJn
vZ5LxJUmHXn0UIH94fNblP2CMHaId84efE+LZBwhbSIKy0CS2B/002EGA7nVgQJCfXrXsJB0NuDl
TwvFklCqb7DvisNJGIR+7H53ZtW6640Lzew3sPdEzmM7uneX1VYVcdZkNUWa4NCUWVLg4udSHGp/
oy4+DrAu6Hcw63bzY22POabqTXpxWT6WMXk4pdjzTQsVHAkoZux+jIFbRJCSrXq3DmHARIDw+cPf
NglPABm2VF8FGUgvbkWZE4lN0JHrHuLizPTC60Irrtt4RHIzuf27eEfqt0hundOU2y5DYnjHBknn
PJON10rU/i0cHil+CkP8yK7QKt3BlggeCXdA9mw09LunueZHiY6NQnqFNYpxnsdLkjykDBWW+ooo
H3V193TTt6UE9kYRgsbkbOGvUAoAVONuz/vwzlf6e/Dyv5/tz6fRpgsCHV56547xGf040FmBEMRl
gp7b5WnSGqvjp9DGkD7CygHDT2MaDWRU2rqE5oye7XtHOG75sJgwbESyCnRaXR+nYZj276wpBoOH
YV4fvX95zSa1+qyvOjso3kWH+X0UOdZDQ6iUxTvTK8Hk1ShDxqJPein4UJqnav94kezT4EJsDzYu
CxFc2G27oGdrCxMCfK2sS2MVqba8pdztLSXuQzRK/lQLOwYMXNaOhKqVnXb6bpqwqEF2DsIsrxZS
dotHrnVudL7KRaP1lhJTV/Vc11H/wLio5l9cHO/YZdvE9lMJLAbmSQnFYRL77qIYAxgVCN9txot2
A0e4gcs2FxIv1oJQTVQDYLxFLxMlUaKhiD8XavHVYzXXOf1MYUDu//zPryboErzRLm/Q07SlAZKF
CfMqBsR771rslo6CKzO3LdgjigOj/QBnEz9m6YgdO1KwPS644Xjn7asBi+tG8uVRf3ltQViI3bDq
Fu0scfjvuC5UHQHuC/SQLtrwu7qIe28RboDMCDF5iLieOMP0WE1pIkW6bGsNwdoxCzKI61XbK/Xr
jd8saLPXY8zEb0c3GiEtVpAQIOhbGzWyBNDV0TYHtY9BndiZ9cikVI5d80t+PwVNmoMM74p0Hkt1
RXKY0MUOqrdOqsdopCKplqjghRY0NLIG+AqoPFc9+SiSLqnWcHkLmUo8gxFzFWRqKjr9ffLL/el+
HzX64KxJTGZLFDHiDFDZtmmWA+NNpf6yIwg9awr0GueDKghuhQKgnyRtltxZO77phKgFWVXVOFmg
p1eWXKf1tFpf+ncNHK7ByzCnGw4vkFI01zVmED3RJnxs/qm453KEUWpa/IZDA3mKftQzGvN1Qh7c
PkL5IwmO2hPvJdcgaK6nL7jnV2MrCerVxp7wR3v3jzD1Cq4A+mKCduD+f3r7EtAfMtpE1SRipe92
MHUlpscLlBKzDVrD4op/IY90x5SPSDbuZb/Lw/nl6BbxzysF+y7Z/YROt4zb72MYDyxPyC9IEzBe
DitL8b1S5KI+9ZJakZgUs3RTvWHv4YMOh/aw981Cje7zn+0X2feEwYMcbj5c9texteTQ8WJyhUQg
Sg6oT8VCxEIip0ijCDVSRTdh9M1B8UAcnOw5IHOgcCMJGTFRv8bktabxmsub3kisz3964tkwJFWq
7bsnCfJ0CRdpLazcURVYS0E+m3Ki2XW4RFHbmdDW38WygQskAK86PVCEjthmpbiaeKuvdwEUm2sB
pk+HV1pWnFvwVS+Cgbsks46n7Qlsur589WHxrJNQZnlxgxr4nGpal0hwaWiwjScSc+bSSBk4qAVN
BJkHpcdkYPOom30PDTFkfgYXPxl89sSds1v79TXgfbW06UHVKVmO6TH2Cpcg//WGk1Yj15uuLAGD
JQ7CUFmiCVZDgiDMY2lFFiEllo6Z7RSVLUFKqmUmRyV2UanXTKzS8xVUFiagkd8WD4dJEF3pSDDV
fyIkgrsFFXsRffBnXX/TjZEJJsaO4GZxxxTr64JF0hNQRHk6IYulhB9Ta/4FqW9A5bDHlMF6DWu1
XlZRIqToz+N6eSlreMe8EnGGH2r63DknmstKq3XOKpfQIY2OwMjRwB/qAkWnbKvHXkKUXu/iXG4I
ldcK0dhjEtpvmm8oRICLG6IRF0qjRyR28OzEZmBJ63gZRPu/buWg5xg2O4S/nn/XE9w6IpBpTWD3
pxhBGWwdm8oAkjp9cMl2F7UqCkwmJPdUKY3Q6lFt86FCRUfy6/7s2mw96FLNJwGC1dK8DcBdMXfT
SSfGT9Kd53YdukwUFm5ZdIAXY67rPXEEgKgxbjXobfAJOBymy+lCUzRI4GKkWEwvesPTJxh6HsAh
elgSjbbh/RhHxYi5Bv/K3zGFheauHuFTL4gbXeFUsA6Tlc3dBRv0Z2rFVB6XtGuoRZJ6P4BXl6Tn
mx8B9WwVVg/ueTZesL/1ggyAc9JL2S96jzkbAFb93hSdktDw5Y8YvWRaugJjqNS3ahPWf/fjZEiF
QmCb0u1RJvUTvYwUVYnNd8y67kna0NdSFUNMnrXj14kol0OwatKijj0YfJn+9W+X8vV4daZg+ZAv
bp1azTLprWsgZo5tHwoMbMBJfurFMsxRihcLA/tLH/nDOh4hbziXndunQi7W6YrHCx11rZfJpjMJ
1gNBhtcUAsDw6QAryKUWnsbVRCgVsMVQ4+bYzJe5UP+j7ZF6bZ+2T0kCspHjNLbWDxwINFjxnBIw
uzAla6XpWv9xhUkW3bwe8s8/q1pH429sdMH/HecUmvze5DHZlwpPi2vSTDULo16QuSNUMNzzaFZt
QB6ng/am7rc9rd4XUIcZ3EritbgOzOEsBkYNdNI1TjvmY6DTe4lNf/J9+fT9kuZPOtY4+lbo67sM
3oVRmmYqmHXS+hmbW4Z9v+IKE3STPqNI4iPVFr9fSumYfpkErJdrX2SgWB03ivPFYL1o0aNxVpul
qsOvKaZrTvbeBKtQj0m34gxHTuOFx3UPDaZ1tI8dG9hvU0B0CkN89Ar0uCvASbM8dpAsFBys/cQK
9oL9oUIT/uMLPIJxbqaYpAxVsfmhOwFBV3Cit2p6fibAIdVRZSoAyP4IzZDw+2fZtPbYJcwwG5ZH
Nd5mOmn/cY0Nn7xFCVa+4XhCsiM6J9p2/E9er+C+d51jOGevnZNfLI/zcF5+3J1RxTuoP7zb8EH2
IyYnD4f972tqBPBkDHAjX2+a8nBDaUvlauChat6Jnu9wFHh8uQZQug297Rsv4GGXv8eM3yLdTs+4
Q097tQba+UhjjRgV8nK42VlCbGkpaPx8VcBoKI7vo/H4wBclzrwAadDu1Ei/4uz6SZBQmC2wcHIj
UpGCXKd1m//K1qXumuJjauiS8aY01oTRWdxzmcB2GVFL5qoLqXeiXXnWoWtfCO6bp2yG4YQ8N6wG
UK/MM9INuiQGj268lzWofxn6PGRyY3jprIxzXx4KbjkehNNTnXASW+9UtYIJL89uCZK4DsLwcDsD
9v3oCCfik/WzG9Di3FvEwdW6L94h8lLgoDCV7wiQSS8CfS8nUqya8Zg0kCbJKZn1NHP4R7Ibhm/n
HpB7N/kH0vo9IKt3G++a7kP1KeoRBvuHxSxErazX+TDmXlX4iTM6DGnebWnJ91uz5zO2/fEDMLjD
eGr+Uxu67wj7WgXc5H58CEAT+tgZKELfqAWLwBMaoTuuNDEcSTnA7x7du2ePX0Jqaj3zL2+zcc5j
vmMfngSRflHYUv+DMI8EkGqm12OJJhCeSHae2AbTnBcbEMfpTAWLUBUMgxBVIQteffLOyvrmXYm3
MvC7OPRTL92Wj91IAGYRQahmcSffj5o41EnYF5cAHzlh04BbuKu9ehYf7NzVMhpLkdAlpbHRMZ8u
4D7BZd+4FiZvIE9as4jGjYy2M9fbONy5QgtH/Q2BgLEb23W4wnjl5AFfmU3p/NtA+OA/VoPyW2cw
qV5s4YCzFHT7uOT639Q71g8LtkmpV9VD++G+e1I0BNOWHIPHDBMRpyvQw/hsAzYiCYY1doIyW9Ca
9yzBafSL0fK4vbYM39gOGdgvhJgfBQTFDIJjOFcwgVpgo/5lIMgUeP5BKsqG5pWH9duYiS7f1hK8
NZhxygktZT4ZJDI4IEqGVjhj43B4So3klfK53R1PmLe/OWqvwsCIJJ2y2M+qLKfwpgOYHCywYjeZ
OMGz2znqED+N74WGDRAKAi4j4ehNyUxlOBqCKOCGaX1eKkpuluMUlHX/SWpAOybdD/HbOL6s+BI6
9LTLv9FRMWox8PmWSIa/E5itXpBFyHN0MpQyw9q/4V32cF5XPHHU5X+nVLFpqiy0J1Rrc9aYTpxh
qaA59v+F0tkXe8BLWYL2Isj67gpXo/GZPanb7Zm2V+SGGdwqSKXbFC+fjeIxII5C5vmbsnp1Ho7m
sWUKWs+OexxylpruXqiVlBdTxKd90Z+8Kjw2LQ+jwtkBAlUrUrOLkXTtAg9WhG9nnRgGDYlFo8EE
wcz2LtuayzprCp5OGVrVgt9i3AGyeQ5MATEY7BfqS5L/ghvIvaZGM4zS+zIegDQsfRfMQlzHIbYl
ppEenckDKJ+rDFosJ9x86msf4dTkvSaajwwatSLrLThB9w94GOA+2TN5GjalHaDY6xfFLobR7Lrt
1RLt20+4md3MCh/7v3wtvbq8uWvdRbeEQtrPVWUZlYDkQM6bWaPK/VggGpj3mG1/22S8AQ/YZeSW
cx5PKuqJ1ZgTkisF7b3AWfq4gyJhU+JHJkSImlsZxkadveqALjwZUMvt03b1jaDcT0fFs2zhqbtP
kbs3tl/dVmqE5au3iuSyusW1Ufqb99R7sUbKGCK5Qc7Ri/Jg7M3PGqI6K2unYnCeL6ccp0J1ahGH
BHjUGVnk6GrVRvvOm1Zn5I+/SPqTau5pXn7Ql0SITcKXqOLUiX9dwOdMi8L1ZuUHB58vZ5SuXOr/
FcdK1F/kVHLSEjV5pdSm6PMt92kjUioeUSqsT72DyNu/Ev5bTxCt+K4YzLJqO+xv44hplNvuKqDU
1abuMmsYMNGYM0Ga30J+xwyKJLfy4PjuIVSOFv4loaXZisRD1J7bU2UNSUUB4e99MkAfJXj2a2Hn
9+lkLmt7/1F343p1odLU08XJ8JrRuJcDvti2Tnk73nCn0ep8/aV6FAxO4+27VtaB1fL4X1G9kFjY
X7HrEK9ePA4fgEL0zsHBskvIgDCPZK4p8REzcQwmp4ElOcbPeZg+2X3XTDGavSqqQkbfKUu4SNJr
RyYc9yaT5VVOtIWZYHb2Bjq7g/Y7hw3bqDoXPGClpCD6/XqiVcwWVXqyKfNO7ikz9icnhzZZGs5k
7PjSw3+kEGvszr3v6cGdtkvcV1dnNe9dq3/uL2KJwz7mc7e1hf/fKZ23jIqO6crPsjEwZc90SoIh
R/xPSws8GRW4UAFwrvNaDc1NDNpVsybjG9bveOb+f1twZYVkDDc4LnMoNWAswaw0abdXrEMzOtdD
neYQmlDZFo6nNvLHRjcdPgDxD4J9HskxnzQxaxWG/rpNkwvVIQaDNUULzS7U/vQRa48F942piLZ4
9N0YCmDB1HtiEe6PUncMI5iSupP52eddw6bp0auzxqDzGu48NNKbRoZjyqART86g4/jI9PeXk3Yr
zEqYl/7Sf6stACyyA4SZbprRpQHKDtzs/QrnbiMg19I1EHV9Z87zhKQ3bf/MDEhjKo9p0elmzdPf
NvClryGhlXDJjt9YirUvmUf14ey4qMCB16I/ESJ8tMpR2wDZqFHw33JspI+/+WzFaKpYpTGS9bub
g5xtmD1SkHRi8B/Um+GIo39wR7h4I2hTT7D814m0+gK40Xg6eGk22mbB/bfdbNo7DqbV6ChUgcny
jzw53RD5bo10FYCzqQ6tvfASSZIz5oQBaOp1Kj/agIbbMfv9Yl+4rWoJn2BFwCloQHMmXPkx4NK+
Ipu76m8+nSEmSn7btuevZWXRUWAnCZrBppyhTqEfKwy1H7UaiNrcFK4Db9dD+OQbm6VmlpQcFrtm
JisRZXCYtglLNF9U6VNnkpnlpcdJ6+bnoRE+K1Ddxwup4o7Ro9VPl5BoW0VjI1G2Z4SNddgIcepA
owcJrdK2fiWrvD2Ha24bzehoW0LT27VE2S51DA4ARPR7qUozQXGDrt4qMvJXqDbXhjeMYvIYCCvt
EBgNnjYzpgkwbnpNi7j/DdoUA4+3Py3An8CPMl7tTKZwm224clpoTSp5incumZbdxyq9itqjL98F
ZQYY6/H8fOF9BWnsLsGvgRJRCjFWSuqy8xS9PlCQUL2T7ZCQV1R/Wj83TmuzjS5Zf0VLvVJ8JAFL
w1m02t3UAF1u58gX8yC2W0lJHCc2GF4CcwREybSTXUYI0SaFXftSpMmb5NTzuErL9CC1ofJZyjL8
d+PLJ+npMrDWqK1K59FS1IS3KSKnyPbpv5Icv0zaFY2XTUE/m9sL7iU+FLlJ9t2Bk6EEBfQZqKS8
82xXS9V448I/9kUcD91KFxFSVBHteZsPMxQQflv41YzXIF7aN3tyaM+5XifeFQ4zrDMMT0NlxoPA
JHRMvkPgXzu+3FXOdIMhpIJQ/DHeLerr5FTfmsOHj4gfpchrCGiuJAKu0l3mtGXHqV0ui/zT7jVs
CD/aI5KYX3m+K/4QkwnYarsJq9sBSZTzqDmxnJTW2SwixrNSjG+gP5tfCzhr1X+mLgqFBN2IarP6
JZFwbfkzkTK+OXUtjkKtU40JYXE2GDeQRpvkp+aCr3igUU9tf3/LAOl4Scv5AC0t9E3okMv/ItMU
2k1dH6MNOC9herltg7I3DEiEBi+qszedHAnCNmm90uiPKPRqdJGI2NtirPDm5LoM5e4fXc424Uy/
5P6VMSfR4EskM23gIKNf5jP0cH9ocpRa7MFrkq+5LybpV9yS0oxPd2OX/Ik05Aq1ph4xwQDFzUyr
FoBVV5+vRVIeV6EMmbGRf67npBJ3DfRv+BJhLypdiVP7QvwBThYb5g8t0UmO7Vtcg8pnn5Wn0dA2
z3X/40wam2pYi+eUCTRBzB9IMspszmR4GoYYd0bmP22s+6cvFVyV239GjBcyNOZsGN4ewzgrD7jE
VlA8GjqaNj/bG1/XO+7IwoTx2UqdE/IK9JvkfqxL1nxFpHyac/vNjTKLvnoIYp+EB6UKbVhWTAUT
xZfomukjXSi7g4RI6NlrqhfveOxknfTl5B2r2g4aCd4FwJvKxmDbcagNR7qorgYKZSElGSJBlSKO
Isp3Hoz/Xzqro+K8qJvd5gH3jY4xH/zC/9+jI3wjHv26zs2YcXTexmPtPwYj5RsLRauk5WFCgxfQ
uNlk2T8g4btC83jngwiv+kZihLVS23Lfx1OXBC1jiFUBfBXxk71+RmRRoqMuCkE2ZHfmPGldim9+
jq8Ru2fXze9xuZIu+tIeOnBmWamReRLaYscw+kBJXJTMdzBUbN+AHhnMuB6cbFq+hN/1K5+XZwRg
pB8GNabAEGjHNuaawwZpjKc16YRgGJSO4pqWsoDSWuq+Mpedf/p1UXi89adM+ggLmTTyFHWaIRJs
/HMX/XIOcLLe85Z+uz7tnqkioXBoHtZG863Wm1+wdedMj7vnIz1bEnXbzloyCHfqWCV63YRII1vW
aCX1MuBP1TFUqop7iR+Hs4+3KJftKzyuO5R6pZgmVUESsZ67M9oJI3xhGFheCe6RyF2ZF+Gzo6Qy
zZ/E21GqfWkwqCUlMA4LGUz3iyqC+t+ffe45p+Z7gfMlu53Z4tVsTb5YFKP7GuRUT5Aw5+fAGFJZ
p1xke6P28H6oJB9Jg58BgbKqXn0wIHPzbmEGIEIbRMJAJZbXnn7PiVwiCCOOQDveZ6QIygGE7TTE
Z7HP2iSR/5b9WdNue+UK4BJ/7xy7ZvPSAGO1rOkCQrRwn8JLTJyWt1KoNZqiE4HBO+HNUhNbTPee
Df4dRpAFK8i1rXAC0TVTCECIJHVNaepNx7x60O7/KvV6tJP+HBhDeB9j8FAsYubCv7dXUja3Ml+M
BKvyzWOKSaw8Aun0Qp/dvwCva5haawg9alKdn4MVcSMX8hVT12l1wT/J19z47PkPfZvsbfvY/m+7
t8nY2UlgzY0snO0bhQuy/gEY9uQFXbT1XBb2giJahQKz3qz0Gv4GbLzNwJMPFhYeLNC/IpmrqqaS
b5ipv2Bso3p0cIWHHExSKTivQVnNML3bP5EtCADNx2BzcnNnInjk71ICa9ipz8AAv+KHCwqOqBes
3LJF3ewoM/a837iHi6lDZyWQ0Ud98b4Ym2oEf38H6vaGXwfNPORrlDl+wtooeUMfCrqD3Ko1EDOz
PqYuUc1274svsNZZGTQMad1FHSSXRxtsT0o9UkK9RGLqicEgMVlMczvUDvdLfQ9BVZ1KPXeJ0h1G
SOCwIqrpu78Nkg7Eb+LAstqKDFIP8CIdGjLbOwF+tbRCFKZa8sxdQSC72hyc8u6W7qVdTZFW/4aQ
idLPRuIlJH373G3rlw4KDwtNfBBZKnrXDvrptTgl3hxhWXHs26hMi04Tqt0bB/SUGsNFhPt6PQsD
Q0ELO4MoqElNRUzVIaagdlDRcALAJHAxiKfZXoft5LdMyCpk83/4nLVPCfzU1HjQbOjoVRkOZ/mS
EaogA+layZ8bYLdO+ieE1LVYWLLSx5M+PsQXXJ6dY+COAyJhyEMG1luABpVI2j2PAS2GVTnFf4Va
8ASQTCiq+6BFoOM17SbLdnnCZT8L1NeWTgnLeYCsY83iK++ZC/V4aAcFpWHkdWQt9rk8j9MFvcJz
hUOHwKWIe8BbCFIkonuaK7QJP75CyYHuhNQ0bmRELHvDD7PgGdI1QO05nzrUDv2Af40kGD2iDfE4
uzPpOTRlDetyoadEEYH0XwCuFUnVGBEA40Uj7aoMV2evDXYXm41ovb/dQEO2bG2goq4hrxouPCN0
9xbSC37djp9PC0cE03giCHSgctGbeQUsiJty4j5CjH4UHbprnFwCTolRdWwcglk37yH2vUJy5OU7
ZAI402SwrRKWUPK8aJzWBdhwMy3mueVivDER/mHvdSRkOGc5nUh9TEMKGqJMmp4BwiM/MSs5LCPU
XMYexu/j5mq58H5h306f9R5tJ/kHxnIxqxTiEWbfFjpPWWcWIGLWPTTd23YJZQpVzsdO1Av1aKB5
2VrSTk6BaC2Y8IjMooVdlzaf2Ug5zX68EMUMhlAyafcAGldmmulNFEghOLWENX4UG8rnYaaY3dWX
K2Ntd4ZofMc2K7ieDEURkvyRasNxeXU4A/0tZ5LWAdAWwahptPLD+qvHHjUlxemqX2U/oOtTxltm
83kipBT2oum0DpVp6HfRlaeT3Ck9IXogIMMtAjIU8QNN5lvSnNvYYM7tHlSjRb7KYOda0uHQ/yXh
NK54VsfHpRyzqUg75fpbt+mfvZ88gUfPCvESZFW5IkorRtx6YFX7nstkJMW2jxOpVhJywelN4wgY
R36GYTfVRRjxCKGKVyztca0s95wWaV4aez+m8agBLNqQA4Vx9pKmUZSUbxRF3mar8YsqPowpt2G8
8BpGaqVClDtATdlfe8QY/RgYu65XPPQRcHwfwBM0md/ke7YH6NRnH+YYvipMxq11wUQgEPU7oQvX
Rx9zJWD3ZuTsCY56XwI7FxLk/SXXQ1DCTC1DRlk6lhameiAwKtV92mTvpN3/SZyCa3fA8NDbUhgx
K/gFBG65DNWRjzEZeUpx+gOxY8wnIRt7WP22p/SwHabXiE4GRiMKERSmjZw6FaNhGdGIZApnQ+p+
lnBUyR//NsmXaWgyFtErB+uTTMDdyP9kup1srEUMLxzdyMG9Rx65hFypY/jRV5/v2tNk2oPc2lzC
u629dVmdZcQ6YnC8ITUte/j184pa4bwCF7BaUj0dK9l5RkoahHl5qHjTA4qZDk6gZlmO/BUlCTZd
EmWL0UITde2sCIHZ0BRyuNCXY7EEk6hCJC/ZOS5KLbxHKzXg9sK8Of2Qir4aZ9OL7o5DTw92H8VI
hRYF9pO1xxVQXEAmeyePynBAgr6aG1rZyuDJxSw5fn/59Lp4/8Mb/PPyFyI5m4hcEOhZJ4ydppnu
xZaaAJyps9FhpQYnFDBab+KjhHSWCuC1WWuS7gNnzASoo6l1E3QhdVVldhNPAwyVTFFtiDvfqptm
mTv/cuwNTZUnnhyIaILMSHD73jLCvS1dtGi5hWaK4WpU3fZMt1C/f/3kpBA3gSyHRuOYMTi1Bvwh
kOFHB8SrKhsdU7xBTmeEGUJZhhDTVOh5qcsSpp0B/elsgXwtWQCMgkQI/rYCyjDMP1m1VIGxfxxK
GmTJOPmOZLPwD3tThCMMWEeZCh+dXmGYSN3BtyHqluqSoodlhm8sWF/s1JxvG1b1OIcClyvO4Hkf
9UcbmUSt+yo0YYhJZ37pppqPWHU5G+d7Eu6VF49V5pgXFpGtEw3XvNwLa/26q1dnb8ZcG6KjwGUc
hdp6LA5LqDT69NQ02/uw+ZHXoGCr6zSEUoE/eXiEAhmb54/i5NMPCcajPmmWJboiP88ZIASup/wG
K6ngDQ0C2RP06aktQfoiAt8ti79j2XR+TXoNh84BMwlGbX6VKvHO3oeANZWefWJpIA/D8ZrDwmAb
tgDWuJmrSabJTqukUCKlAKmo9VyLuyyFgCsum0RRt5LzQgoaIZzcwtXiKKbuASMt3kkX6UOHBYTs
s3QO2ILwrrSsyIGHNxq2Ob6fcNqkIJRT0wdYrytw2UIfk8CqakNMv3iWl4t+/ke/vXa4nPiaCIIm
aoMLZtpVbCdfPc+DG7HRjgvMy0pNXQC34LegTVe+3Ka5Iu+xAXHgMWJl/IH2faALYodR95Ni3zAk
zX17p9oUiSWprDLliqOwBbMyYf7F2qL5PUZw3R4pjivB+yeZgHTYxlYaSGCJoZEyyGnSpcnoYGWF
1OvhhB0ymYEpG0WlSgU71WAkkpMyB8F2MwuSXjt5mFF1ye4MIGxabuyMyX03Oc3WZKv93iIr1LdJ
JVcXG5lc/a68ecrFJN6J2KZx+CiDyfFCAZn/+mpy3Y/CYYdqagPF9XmxFc88aqRKYjWeylCbrj4q
CiCitD7JnVo0+HVbZtN/vdDAT7Z2jS+XCuLlMMzkmnchYrfZeviBjUpLfcQ3crmpHv9+9PpSrj2u
7QhDhVucvoY1n7UvPsTz54jEyL1yU//5lSmaDdjBmfwfpWlQaGCqHZuEKQefPr59VN9uiJ7eRVcL
N0bkjigaPZ+4YNgHWsvRrMPDXY59ZTR+aDd/NCuXlMZvVqL7OoEd5oYvjY1UwHEzXGAGrbRM5YZS
Wo/fma+2a595bZHGkkfAezxMBrF4YRlaliuRYFZ6inBfG2zjoctwoJfZKMkDGoud+qAZfTS31hpD
8BqPmhKTYphjYBJSOxWD76MCVhKplQjxJJFZjnRYhDyzsIJfs+bVPs0Tj97WWN57fQRXDeuWwFDc
E9fVHUWve/V241NtVg/LlKselk7n4wSd4d1C9JZb6VHP4MMRAjIPjzHmVGXUh78xP+TFjXnBp4s1
1rUZ2lWEpPpb+LgQeLeKIyfKaAef6WvqGljdlST4XLrQUmP/TvBspyjJoQJE2fsXXeMnJhAv5HA7
nqbz+3gThlEbUZXnMJ70CweyBtMVs4SSgioSkFZOKOGDAYdYc7g+6cy9M4pyLJK8NP6orBXv4jML
0tCYVZc2ONULSxBseIoFj0hdDcGmhYhsoPAD6sxW+4h2tJ/E2nsQlxgFgO7dwCOldMOBHMGsZi4R
alv1Yto58Rmidj04q1ouPq1FY+h8BDnkc1RYncQsvXcM3jknWTSI1B+/xNK+Ie2xA9U5yz9mgkhs
AUjtgWKhpvJ438rKsf7ndXVCzIzBJcI4CwII6MKYIzK21z/yeETE3RKRFj6KhL2AtNQjgrO0+mXj
heWwDLw/xvvdnc5YHN+U8YcSZqu6DMujllESuOn1PMDNxklZwHrGnRM/R0+Z2Q6uDXenvsX9SqNY
2mx1cljSpV5XNBULTMNNc03SRM4ZkHkNXP2V3gsE6Tul/xhIN0bn9d13a5kKFGCHGoUENg4nWV0R
qzHY7L3rnvQR1bBzW/oDczH3RzizZ7Ywp859CgNAnfNbCxQ3WTe0MEz1/ZXcZN4A3fxjM3w/4oVT
7mUEhumWCqptyvQxaQM6WvZITQ8kiPM7Kf7kYQwhx58FsWTtf45to2aUyvLZJRJ6IfuAO4Nx3Do5
+qLSFmZqTcu+tBrr+4NFHok91extzyrUKN261v+ViHUsSTmqB1v8sySprWffL/Og8zznoCIWMvAZ
/RHTwVPLykPzZZkoWoJNmwH57yacyfXAUMZJ0c4VkxlyYDkUy+ZMTGmqiYBGCC+CI5I7iUC6giUE
SQByDmdNlYW+RZYNASRLmBKOjBjdM/zc86OtgqlXC2rqMjhFaZseT/2wQkdx3zVgqNT/Ui8krFEt
C3GgRoe0rWB6fR9MYSHTuMSaVbAIt2bU5xISsWKNEeQphXEcjUBV4NcQwLYYXj2pIkDhjkRPueQV
LQz2xeSE7CGQj5OVvSLVQIJfnKfA3ji3h6s687UYhv4jcD44GwPsaZbAQsHrR+Q1u9IkdDx7sVXU
H9kz2VHfXo7InbvLDScsYEH+/ZzzLc5EEHQdlRx8C+7K87dUVl8hLH8mUHy48R3LFUoaM6X9XKlu
ti5dboyKx6jVIvo6/khs0o3Vb9P9tW0y272K5eU0490yg42UbZC+xxHzSY1Uj+sAv60hXEg5nQb5
o5yjZEt2cCFqppEiOD4jHWKXe4VDK4iFwYBZ+GRTrtTLn0h0jKTyM+eLwE/tqfMZobh/ZU5NiiRE
+ahZeeq9e50oEEPGIX3y1J2qOu84ZUBgtnaHpCRJTuT48aZ1K5aKqGlhZVXUk339RQsgql/YFoYf
vx8xB8x0URpcP1PPbESGQA3/5RQtjo2sax46I/K9LKaeQBln1X7ZJ08mOWsTBHCiYsNb6/MJrv0O
xILn9hS6lR0MmzZqdHl84phmrIi55OgitW+ZZUaruXYgsPKIu0PYmyjnoqB/kHOYBoX4RKF1ZFOz
XFd9N4hIOR8nb7z6AMBiQQ1VxvCK5M71AFmYUYyHn5v9fpkQWFQuY07H51/deMF6IrsLYPFOfQag
yN7BXQdBV6vuNLxBAlTdzMFKJ9Eb/wf71yrODR2ezWsCDPtOp9HBb6df1+Cek2on5WSIH6RihGeA
eV86UL3Rx3qOZ/5EaRkFQbYctZsUhwoOZQAnYZJMsBrlosomd76D9Q0Y4jiwan9EZQLduzclWWcQ
jk9SqN/BzdtjEuMkkjXsWlYUsESB23jEsfN5IDK9xcQpae8PcuOJQAePFAGw8BQtqE4wso2emmbQ
ibRsrlUaVKYx2yVOfzkChx8zmLW+NYBR6B8OTBaqLQKuVXL/r8bOUoecUB1MjEOIuge5RT1sQmUZ
cO++yzGkkIqguEsySMfGQCAKBrLVYcHAHSOcyJJ0ChP3ywLPVACNnc7enTFsmuEURM6kyrND3ArV
m0Ypczjr5ms1SkwsSCSte4i+u+G+2coxi5wx52BvINix03AfFEO+c9ggNIejNDkyww5R4grK4GYU
2nzrFZSddedhm0P76z2TZxtFnlohEOeIOfJ9OvgGFV9e4wgrc8lz51TTCFqBkpg/BHzG+VGYFs7L
B5BrmVKNUNjKcQhHWmnf49xSDRBX3TjT2RPCkq7rgDBzDk1qIsyP7r8dQb2+lJQMHI3KMgHgN4I8
3GCcMr72kMVULE7N4m/ZhOYpU0A0yXU9MEwwMrOWbOrk5Pr9letIKAMWIEo7Zee9DNumte1/j8Nn
kiPe1WzC/aNZWYwlHLzuQX+VU6v3YC3m1zFrzrKp7LUqXdirn1Y7lVyoQMOW7bS7bASHrLsBhaex
IYz2RyqMrIIcj7isA64uWflKvg6AajkW+r5kttqX+Jis77IOXonzHoU8jnIoqu3dtyqp7q7rIR/V
UQeLMtDvx74TH5W8ydSUIL0DxA0p1LN5+O10mvnHPx7KeZtJLVgn02vqOhj8BMvwFl7NpDBVm00Q
vY8Jz6OL1XYoBDMYuhufpW2kAOWpAPV3cN4BmtDXcrkJ8Ic/v6Nc0150JXjRqYgaF75AFMHEtHjM
I3DGbLHxequftCyDBEawoamC/XVPe3Dzz1n1OUPLoo6JhGtHH4oJTAASGyeCU98ry5LT0gRUhSFn
H71zf49MWLduOEcPkaAyyKPPbR5IUR3V8cKyBcLzQTFT/fl99WVEhyJzEGZjsiImdQl9pwOKK72M
u5m74qBqGm0+oSE3L1qtqpQAPfIwiXa3xE64qzI7K1eNd8/ibg3hsLXG7XkXuFxnRQ9W0FSqbhwc
qOqRN7nLDpcggMIeIphzS4xjwLcYALt1Mxp4R2UqJuHJ9e/HLha4dqQCYAFpF54X/gUrLGzMV+xU
HZe6UNZrbdG2Cua4nSvUNZk+t+sd2Hasi3EnpHhJ7x6mMkdXJ2jmWi/b65YrSGW5IxtPHrd12pUu
KqSiGcdj5FGHo2eK7PfKWhshlAfYHdwOXbS6EpBmxkCFsIQzC+4hsAdI+m/XXFydln0fyakG20Yg
NrNOxZT8CXgUEzLtue2aMVCRQBHZTFksHw3CyBFjq/cmFkgC38315Rwqjm92DOBPT2kHmZ6RjIjv
qkmv19ICf+k/TSxSiURRhfq4oUTOxYNnwcOS86/t0EWvSIgSuAFFQaP7EyU7rtil4ZXDmWfRC2xm
2oBYwY2HUNdW4POqGdQ+FB75LpXvVu3cWItE28mqyxGRbBvKhyIwqvWfdqU14onur/LPFUgBACSg
wLFsgF+2HY+qeaH6uSmI/OlXxgQatMtMk4laRE9u6NV3Xmxa+Jxt9oLP+eszo93dPwyz9vDxP+Du
NzZhcp54piCIneDEWW5mcQZJ2JizlFMj8zRue4+6X5M8NFK7YCJ1nP0s80IcYZ+KnzP3qOhQxKbN
o7NXo7yZ3s/17uq3yQ7+eteMbY2ZbIoxgvXhCFtId8EM4FEygisw4ttUH1EfS7JAInH5UlpbXu0D
dF5cc+R0GTHcprEA2rOjJ/egGsPkVN1oFCwEpU6RV37dyijTpVtLNxD6nZgd6qn2ixd4kxqT8JHR
FJ5enoc4EMSH972WYZOGyagI2OtMPd2QlsTnQx+DPVeZEm/KPVbT7DOv2nod15yrEHlzFeoVkewE
9gaA/I+UE2SM4e4hk0+gmWGJlu7SQtnWHNC5uuHj1krJvbRHrgfSR4HhoiWWfLh97/48lINbdvph
kTjFv1uPKeTMWV/3LXjaDRV/xlQE40DlzlQc6T6K9PiLj5zB5XeOERwFBiNtQMERNUD2RN1Y9eCU
IP5/x1h6Ajl8xngDB96az97Sy0gH9HQZkH2QSTaqJMASNgu0QZPX1bqA3Up7ourbQli3ZWDAISZV
q3oOP2wcQu7frpnbU9pgmdxRv6FxuzwgSPPkz/j9FrNc9+iFwOO6XwngbvII4wIHGX43xismxwQF
cf4JCs5NYQYjdXUr8o96ofA4XKNFBHf+vKDQhmY/5YK76GlNXTQWULSNUa2gDjyGoQIl9at57I43
NeES/zXbSe5ArttmhBJ62uPpWowu1EJkRKUga+MuwuXwYR4E548BHZubUEy/EWSTG8Iu7zhjYfk7
HFigJr/ZvqR4Lmim5Wr2yfgtyXdVkuzNqBMCzBZ+dIVQig/Xux1d5LxYoQUw7pO1P5wxhSNfHB7x
fGpYkUoLrjhrLJnC12Gkfm6QJmFGyz8OuB/wC0Z7IGged8yDtRHNxgvZRRxCrLat5SxfLxsN6+/T
p38j22vk9xGlftZjv1NLLKXQc0dcnr/8Ee3t0QDXzqrvU56R+BHbAoLTsAxg3M/hBvDW1qlJq7Y4
11hcDT6Jm0HQ6UhVzuBmmJ+jhksLz2353OBNy4TmRa28AonUxl6++JXuyCfdSEpsFjNuClIJEL+m
vUbJmyrmOJDW4mpZRQdFMqQg7KOETOV+Z7sJMTMfI3FlemYBZjPZNCFcg7j2N77DHGLTSAei5VPy
4qyCyhl4Wp+b39R4uEan32lACE3+v6giqIEGo65u6X0WaByDrcOFOPrgGBZAlh2cBexLhs/t3ZYm
pkeckYN4nhfjkFa0gEbuR2BMbiEx6iZqnsJE0JKLAtuvXjDfO4Nha6IhzS3gFxk5lSOO8luMdhRL
C+moenaufLV0lICOhbdu3NQDYpw9wEMWhIJRyVg9qnsE8ZAZ1xkxdyxgdhMku0Vqy6tEN2Eon+3r
cQphpyE/Ji65wqXxEworSH4zuZ7peeHcGJmhH5KS3hoCy8EBdMFLQj2VI4EZvgikF3jCOk4co6cH
XSMvIClfaZBZH46P2i5/HEXNb5NoKwjSZw7d+aGpMX/xujRitQ4qHdZhlrgJ8HfH6B0s7XqQ6AHR
+y9DRmh2VsgJW+oIj4PX/LPagl8MUxzj/JVJ0FMIJV75XQFrG6D7fChilQ+UFnDYrrqsJhOqvliP
nXb2migNdz89bPQ9jGGeHXxqwvSjArXl1w3g093H12IFqudlloWacUd6DowNu8RHDUp/l+m1xEkh
qQEAk3VdWeI+K2ZZT8gAhfnLQ9Pv9cJgzw123wrmAso0KJQIykUmaiRw/bMx3NvVXR+SFjpO2bqs
v1GBKIQC3VSQCQM7tmkS1OpYLv1GQo6C5/d1YEYXo3TO3b2F+phUj9q0VW331oJoCUTIDBc7I+Zj
OfAJwtJZdxa7Wa+iDiBcsyiNODNQxxmwXzzodq+xcLSUtHVtSyVLlrUx21ULcZDdsOEAtU+HWRG/
ARoenY9Msp3BdP9C+q8SLK4W54qEOQmSHQvWLp78K/75YH8k3LypS86Ja+Gk7Bl82/BxtaWGSn8q
d/J5+6AABtDZLZ37E2MT0EJXsOgq7TEfoT+xTGEN/+JH0ySnqJKLWf/gu53nkyqV50OB8xkcaBus
nphe1lXOC2wNh7oTOOB8eHG05DnGDag9FeJsI8rkC3DOfR1J0131exl3zjdd/n4H4Nt2dyUUeht0
MXl78ADUjzx8Hi9NWluhb72BUA2iRh9Zonb+CWxdxuTkgcKNS8vSo0y1NEMTV3zvCPtjF2Jzt8/t
3os9Y3RFAM+D79/AVBKZOx4T/SSGc0/USaabeEMGntFf+wVlumCRTrfaGiSjLE/jAVUZgzsatN+Z
cYIRqGjWGvQmJpM5WKM03hMGACdKz214ioUKjg6waQWwOdeaRLEajp59eOTogpGlvHiYoE26L7MQ
DYCi8h/cbjzyGihwbSvplyoi8jsc+ZxSORBKSsAr2frI4bzA8C7/Ea+iTr9/mOoXYgA25B3rQpq1
PSGggu+Wtc4x7+SYsDpBVLLtSvOfdAu0xBnEEsY3yhSzoPtPplJHt5pupfVA2+/GF4ug+IwCpOgj
Zei/mVDMsULdPAHnwtyuKq1DdDjIAC/eXPOCr1hZDJylhQk2fxxImleE8fhYe4SIwAjy/9lt39OG
MwhZPKPQef69N9RJ3/kf9AHdKwsPDc4uosPK40l9MaI6JO2FBzbobMBqaQ/l47trVL7bJyxiyb70
HpTKVeRQ2YwBGHTg5c/09DngOTQ4Nd60+psKglbIJ2kT9pyZGFdEZ+nb14azd35qtCTCsXXBHtmf
CrP69iTtA+EXxsnf809dh+k5zZW0I4NiTeOOapQoIYOeel3WJPWPOjKaVDHfM5x0JgxRNozVwix7
fGxz5jZsgHNO0+6EeIz9gH0tYnzsiEM8O2aTLsWPlF4GLKSR9P1+VRUwqSTEaqbVnGAxAjr9sfMm
+fG2K8u7/2BkObxcToDChDF+eNqBSJK34En0W0fy9GRaNVkLmY0haE6QfjZwiFQGOCFOEM88dBjG
JZ6CjZ0cmNWKTIez8jn/zbdASzZxpI2je4NypaVqzbHxJeY+ivMHRq4Sv3mN4cPmn82XbYeqa0yV
jeEUfbHuqr3AriWQat0B0y0q2/9z7Jy8J4KCmFdJzFyPRL9hzwOE+NoxvxfzgKVSU5Cq7JOmLA6Q
Vsbx1MlDTGwLgH4DDkzOQFySduYHfoOl83cS3X0ytCdDRX3pRua6b64LFaFYce4L2L74HXRnPJhC
L1/BOyTKir4Z5nofNYOAdhC0i4gkDo0ADCdKFiMBizglhfsLmG1QiUvom19c8CMYsegp/Flex8eY
nsetPSx3Jxvjb5BxF6zw4KdWBIRr/ON+avdJhb6VHSyRhSbX8U5gIui34qXdC5u0wTSbu1b9EiU/
oukAEkl+T25DFig4HejDeddaCBtwUSQQVOA3PXfCJ92UUyoPs7Mj+mpyUBLWkoh5ITZ15761tdC5
QqHveM2dL3/CPLw0p+chl0lsZ4O2C92V1XR9OsSGZ/RBvAw5s4zI+kdkgu4m3YAqmXF9CVjRhlQH
Cl5nxE9HPF8XxPtjw4HDwSxj8WDrJTOAjN4VrMf28C0RzCMzaE1RkejQh9UvVQoN6Bw9t9jQUzua
1wNmlnq/eFDKO+6cg4EuNjhonqcYaiq087mhBw9Pr+Uf7CQeNJ6ZbEx12fuOx/GafAMvOFSPmZWf
G98Eb+YcSVbbC7A0gsRERJzAR3fXlFm5swgXbT8i010GzN4BxD9BVEkLy1EQADH3VRB5VmnXDiUB
DSA0NDDF6Eds96CuCVPQPcexok9+2Vg663UhL6zLAiAopGnCMxmqzLqXlCeQppOI+0Li+OqdbhDI
xUk+EnYvOANnboYYjICOx3ywGwA/+B67I/iguJRu+8N6GFtO4t/AsKf4EhUcCOlkekdPp0KH5/2w
4DKN9g48P8aZx98z2m7tvgt3uzLix1chUbCzfHFIyzu4SBNLujSdZBC6oKSGEPjL8p7qxVEWOGst
Z3ou4ygwK69vrjE44TKa0Q3ADA/jPV9tY+0WRouYNWaX82OrMAtkmbdlTaGX9ucHHSqH1ZJHv1yz
tgwtptAg1+mms5LRYEnfVAgNRV5SNcAPGu8jMHgquZqcEiUOd8ftrHr3Cb8R38hygjtoqEkPaKUR
iW8mkkIS6h2LIYcXdlYKvu3s0TPS1RBUrc8jHo50VwbfJohl2RxTy7mE4S7ovYxyznO5yEV1nHCV
sOZaAJfO9iYgelsHi40AbJNJSs7Wd0BfmuoL3Vonucf2HH3SPEZwFIkRL2pMYutJl/f8twJWUMnJ
RTjnbpREPrJ70DqFPwUxNO/CyacfRkndTk+WzaroH0PesRpiRoui0RbtlIlj6Z9q1wq7+b2QZq4D
y+Behqk06J1ga4ZxiYh0OvANVcAWsJXXBu7sdzRvcWsE0RWB6NOkim8875GvcOT09HtGjmtnw/55
YOS1IHrXIzf78GFnBNX09p00InpVuZW2xtJeUHIZbGIR/U2ayF4RFCx7YLB5cOOFpFBEeytr4Jt2
bpVVH++XcXraSMr0hX9JAgIDOmhP20Xeyy/qfW0ePEb5Yv33hEFcG1pE0uAthb0nv5XfvHSM7OPz
cRb7VcmOc7Yv5Hm1jEoeEs3eYOT9qoDNExQU1tb4DOJ/DKBbEXkWPL2frLKOOtbTzWeI60Q1C8br
2311FDV1VLZvjwXXD0CgXhcYs0YEP5klLfTZLNCswTw+Kj/y/FJ1m0563F6LBuVB4qo3U0tg0+Ln
QR8ORgMqKDadlYshVrNrrYL5Yn2kGZz7uMU/wGoqfqrMKmXHVMdt9wXZim9PVEuSLM6dL0aWtnGt
TmKSIarWvA/VRkslRpfwcNH6EoXUUlbcbG3pe+TdUITvIo/g2JpDo51EZV+6qJTkri6M15SKa+rj
Mv6amM9PsPZ/FyP/5SLc0vpOsgAKZlZhoPGnQDUY3svdMKUrIAvHSq3ahkyX+h2F1ByRLSqW1io0
ItTvMPLuG+spDrk1KJkRu5mtAOf0YlljNsWZuQLOhNXoJ3Sd2HDm/yaVlyXJ+GxHEmPWojhLbHpC
XIzLkbb2o59YSRZJQn9v7zvbZ9oWzKb5rDSefYyPn3bBkcGyIFOHd1ktKXYFJJDx+tGYaVbGKP7P
VW129YaXZp5uZQWswDBy1mPYyetcwZ9WKJO9HwCROI7sQaMmS6HCqV9fkFPlVjmS4z85RT7x+W1M
tNqjyfFWhIHSy16ORD9Pi2MeIM6V+p08AYmWmcyywBL+2eVJ832yTA0CKfHVOe6FGyvAh46pmKWu
jsuSzBDbosZCEdye97YaMnYDdBMkDq4V5uTO7ZfnCyDucYMMY8IArb46kFjw3QUoc1CQtpnwcFv9
gj5mdnvye5rBh/yFujXqDzgqMjVzH/eBLdXrMe9ttpw30eHmb75VqczfGelf8eUrQ2PKTh6XNVo/
qc0e6V8QE4pZg2e9PdwRVVVZ5Rr64N4mK17ts6IYwc/MqsQUaPsT7uuAo6YhMDWpNKQ+c2UEoZsB
DMEOd0LSoArbaXPscqmX4raFBC3fLxIT1CoaNW0ag3siJONGfxgC09FGOdUIlgfvCDYAQ28H2GsC
UDHpePb3WgDfF+ZU80H/y7Z3dN/PG0kFZDd/JSRX3H7WBJ6IWpGLwIrgb/1sRD10E7KrCgchT/N0
MXYYBCr0dT2qqG/aFEkdLLzicjWubYtyBOq5eMDuGv7ZEb0t/jml6xNYt3sUCA3aXWOA7mkidiq3
M9Lz2ajCnFIEtN4jjxtUTqNPwAWNQuXlCRj/JW/V+lZbx+K2eNkaVjxG7g9nxJCoiCt+Q8kusfd9
Ea46sNyCTPObT8lKeZX1a/BuSIlr6VZFXkXjr8Mja+uz3GlZ5sf1v6ROoLxiyGP2fssmislBCjKh
ALKg45DZtqlo9v1sNhXeGAIVpOw5WZEFpGh39xThAGRpDunuz36FTU32Fd+Tg5cQrkL7Bwkr2ewr
r9mrGIM72rJMZMRzAkSQ+wieeolg+R6xY6yldmY2t6zTVVST
`protect end_protected
