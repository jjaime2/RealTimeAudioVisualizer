��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ���l�$�'�Z���u��E�a ��B'v/�γݩ%5=F�7z�N?ysV�k�b#!sI[-~�G�m��]v��G��&��qx���m/�H�w��V����f�Զ�vp��B��\6�Ads�-����jfc`�kQ:�k�ɭ�|��&Υ�B��n�R3l=���]�_���Ro���*s0��|Ft�m
D�e4,�t�N.��a�˽�T'�C<`�e����E(�!$r�)��}�����3j3Rċ����7@�(��zmt)�`��L���Ì���j�LWS�g�K=.����xjG���kT���m"ˮ�vq��p���#1�{�=t�N�/(4yG��/�137o���_/0�����g2��<��ٮ6��S�m=r4�)W�C[������\iV0�g��2��WJj�̚����4j��G�p�Nǲ��˯�q4�c���E&�-��hLޱ��h0�@��I��ǇC�.��ΊvvU��������*�pC2���|�*):A��k��î���#�Q�����^��[~i�2Z|8r]�s���~��sD����*&��եlt��a8	�B:)��ٝ�NT���%%g�3Bkq.�^�d�0�]�3O	��bk��R��4����'G�l{��?�%����������Tٳ��ɋ�Iv�8�L�*��#%'-ímC�[n�2f��k�6!�_�fBu�s�z�)22s�0H�� �b�WS��AưJqj�>g���T�a��
B��m��a�ŸҬg��<�=�у�+�nb�=���a:�� =��X{�?w��<U'�ӌ��Ԇ8r������́Eުϥ�A��@I`�p���^�G�թ�P�e�̈́8�f&X� 	*��w<�����jG���.�ڏ-ݦ�|n���{Ӛ����B���Qxvc|i�'���{ѫ�,L  ?E�i}mQ��p6�З��x�㡻�J���n�n��ʦM�S��$�md�(�����z�I8`!z����(�SCk>�ؗ7v�Y����@&��k�m[�MR�]����$�����5��3��R�fǱ�O!��z�6��g|#A��il�z>?�����_HC�ֈu�v[�-�=�Ⓖ�+HCH��6�b��m�����xg�ܴ5�Q�~%��Y�ס�j�|�G�U�Vul�<�y�G��������T�8+!;h3�=�C@��ӭg8AZP�Q��-9�ϩk��#�*�j�n>W�����Yz�� (=bV�Yf���4'{}�2V#XJ���h!O3�]�CzmYC�X8�m����`����h�1�,`WI��;��-TX�>.}A��?F�٫��_Ey��>�Sr����*%����Y��='�f�tU�ơ!�^�y}q����PŦO�ȓ��	��5�irwQr�(rm+�)�K&(� ��3x�?�k%Z��0߮�8��H���f=@��-�E��kT6o�E�!J�ӡ�]����\G*_(��[x�{���h	@��Vd����hY����a��Ƌj�n��s1RN�E'-2�[ǿ&�?>��T��C�	��]rv�43��|A̐ \�%���.g:��|8:T�����������U�T��[u��(�.���.%�RPm�j��L�,��b{�_gw���dG���Kq�$�b�O�t P��'1>��.��@�L�N;����p�y�
��ˠ���%3}�B����⍺:�U��[-�����,���ʑ�K�]��"(Oʯ����S�C�z��o��#�8@�Y)n	cn+UR�W,��aX?
i6R��� W�ET������s�ʹG�mg�~u�UO������7��9���$��ƝZ
�Ts�N�UN. 1����U<ʮ��n��d#u���7��jP�H��>]>X��m��@�SHteF(W��PU�ͮq��$r2V؂Eh*-�������P�������b�8?]c���%���ts3��YG���^��7!��\�徧���r�+����c�PE�p���Nw7əIk���(�BI��,JзT�9U���bS��{�R�w�U�H
;��-}�ãg�	�ϰ@+,������>?Rs}�1��$��Rs��0VFQ�$���"Yc�m�.k�T~�^H�`��<G�5�"�[����^j� ��`4��|a%�磑��49��}LB����x^P�K��k1Q"MT�Ik��&=�����ˁ�ͱ�?��4�>�ދ�7�>�J�m���c"1U�D���荟�{�+x�ҜD���X��DLD� ����Wg���I�z�� � ���oWT��v[�t�T��N��P���K{g8j���o�_.fO	�N�	�I����M��V�M����C7=��O�~F�ϖ ��-���h��g�5n��%�Kl���C�)��$�[op�F���:/���M��fI�� 1��R-���mg�I�tx��]��)�X�u������L5�%n��y�>���E�&��3������8���cS,����l:u��~A��J����J(�/%p��(B^��Rd\,!*FgUu&sz�u�'�3�5�e֧��n;�e�v�8�?@^O��}�2{d�вѡ�Ӂ�[��2���lw�iĳ[Ḵ�O%b��V���uW��-�����S�--�����G�w��3o�T_��@g�o ���Y$&n�_��.�W�T�1��L����.�β@��~<0Y�	�B)��A��U��޹�D�v���Q��a1�	l��	R&�v�"�}�=�3�g
ez]�b�:	����l��\ay�2���^	��E�9U�֥�5� � :���fc��+���_\Zd�v>����XfF���P_���g��_���u��±��{����P��|�=����>��$ߢ>b��b]h��;�>�k�<o�ZLp�ͷ��&USK������P��ˡ����J�`���l,�C�SW-�c�G�7�"o�X���z�;��*�hӬRU��R/h���,��s+�0�~Κ���E) p���xk�KF�sR2��n�Hp-Kޖ��J����r���(��b���C�'����/�o��@�o6r<�P��N; {�\��j��u��^�y5�wBy�uH�9����gJ�;���(�N���'!+O1�9vÌ�nrlKw�{N�����I��]����> �������3k�JW���T�Ij0��X~��>�����7�Г*ߠ�rF2Ⱙ^�E5��(�4��&�"���Q��ݶi�J�)��3A�^�f�7)5��t�;�J�.�NqV�p����V�r�x�u�HsV؟��²��� �އ�iBh�!���m�W��H2�;�QL��j�d̬���Tn喯=K�'Fr��k�s�!G$D+R
���ɼ��|��C��3��ƞ	&.���Z@"�[�(����fv��_��w��_e�3����\o.�1��x^��2�Qj�b�oYI	@^���g��Э��cG�H�GS?̻l~�6������e�p����J٭)^�G�.ɛAFwfl����b;�1��?�o�_��15�C����o	S]�I��!��na�Q�D�.���@���\���2��.���ַ���w���q3FC���ԑn��I=hb�mI�,�s�hܽk{w���U�)���'16�yk�%6�=[em ��#"����(�,��B�����%��Ԛ�,��"��y�UN6�d�����sjI�W�i�;4�`��1n:fv-�*���; �]q�΃9gxKh��Y̑�7�ިAx�J�jPF����e���x?�N<�o�ҷs+%W�$2���d��¬��=|+kh�0�l�1x�5���tbK����q�M����A�y1Ʀr��e4J��$O�I�w0h��T�������9�{�5S-�k�$*[ؽ�/ϐ��<71�I�bU����b&o�j ����:hQS?i�R��aT�m����T�|C�Z|�i:�iSmT�M��>.��Q)�a��&׎B��<i>�����Ѩ���I{��v�t×4�Qٛ���T������\��tZ%�K�^XI��QO=�8K�Pa��J�}soh:�&�jgU�T���y���l.���$�������}H$���D�s�-�.�O}�p��6�rf&���P��۩�?vGQF�|!�����]%�	c�?$^��\����8y�+�vQH���E����B�w=���V�G����{��c�j�x���?�!����Ϭ;#	]�N�T,����]{4ܾns��l��B-��'y;�M�Ws%�޴�S��%q>JY5�F�/�  �8�=�	p����c¢�X:�@>ޜ a��\0�f��PІ�؟/�1I��K�]�'2��#��$_"<��ψ-� ��2�xg���e�Y�̓DO�46�d��&�M��
 u�\9Q�>�R[>U[\�����=Ɲ|@�y�-��m�֘e����W����f���r��~�?�d��H�&ur���{�0��E�Y��kA �y�ǰܦ|#�Y��:\����Q��=r�b��f*��5KN�E�Mt��L�����t?cؚ8�����D�|���t y�q�B��a���x�L���� �!�Φ�u�$�]��CU �����+Bk�R�HG;`ŧ�^;�LX^r"D�`lB8�����?2��$4������8���ˑ��ӱRR������(Q�@�3Q8��g�WN�p#6��+ڶ%���6��6k@R��6���+x}'�"$ݶ6�6�����Cͭ�
���U��.��:����)!g7K�Q��K�w9�oN_��@{�ZB J�\�I����5{+�.ԃ�υ�+��2̠q�eB���W*��8��l&�Us8[x<�@eۆ���� _@��7lus����!�O�%��~�r�v"~FOT��&p��H協�U%@��!
��
4^��'?������WgO:^���%����A�5�\���RX���fF����B-����P�p�O������u����v��X
�Ih]�B����@�Ȓk۾�zJ�`���]���/�&��L��S�#��'�I�#hVÉ���̭V�gRi����_߆��@�G�����!B"|%�� ���/����>%9�B��s�G+�!E[}��X�����5_W�|l�*x�Y�A&q��AzX2��/*U_#k�mk0����l��̾�o� @�I�M�H���Cj�*e�`Oz�FT�ʬ_��֯e�
Z�=&��`�H7<�]��E����"�r���6��Z�[�bf{�2h��>�ߨso��%H�3nt&Z�L��$�����x���w*.^)�m"�!O����w�>��S�/�2:�jRmK�'܂�O�1L�ѿj�@P_��kr�G�z�h�wz6�3�sr���:�2.uM�&�Y��4B ���ֶ�2��T�9.,����Z��hmA�������{_`Ĩ��^����@�:w"��n_%Q�t�Z�X����8d�Mރ��o�6�+�X5����/�</r�I�i#O[��O�`��s�X�P�7�y!G�'H`p�^��Hy,�8��RE��G. d��]_?Ó�E�9�7���[]�K�B_�~e���� a���cY9�dNr���A�3�Q<�lM���M�R���a���tG���Ʉ��v�!�:�:��dW�j��(�24�L_3:"#��ו#0_��x.P?f��Kl�����W���kg&�q푭�0'���x*�)��K
����V��ū;r���H0���<�d��3���HI�<����x�LCi�7�x�3���;�XRxq���$�O9X�W%&�iu�a�@N�_c[eo��.�[�(��M���>ug��Xer� }��KE�EԀ:Wd�*�v,��m�&�٥�Sv�YF�:C��h�܄���R��͠�@� ^�`�19xќ_�/Q��O1�\}��a�Y�{�6��j�)m�n�>�	A6h�7DL� f<����]#�v7W*B¼��hfI�^j��^+\M�F`'��郵f�N9�$>��P!���NA`Xk����:#�bT:p+�K^��}r��!�n|��u��(���s1v`��{�mi�-��M�'u����2;�(sj�aD�ix/t�hþ���������}!E�^�~4�ho'ƫ�`����� �x���w�Ǿ��aA��)�E��1��V�|Z`�����fb�{S<�9T���qR.W��h�,�/![��/T]�P����W/�@<�)i G�g��J�
�c"���.�7������.��|!	ows[�9&ϝ�n�Uɸ�G��j�mی6|g�����<vhS�L�s��bW�xo5ݐRn�i��xS%P�/K�|_�������v{���H0���`m�ґEՁ;��XZ��O�{ݺ=VGq;m��+��;������T<��P"��q!� _���e�n��A�_^a���
Ւ�]I�EA֛{v#���%�R�
!\�,�ݠ��5X���%��*���+	|���uYmq���&@PY�j�΀�W����Φ�Z�eÍ�׳^(��]QJ�R�g� ]����� ΕsfB�������0@;����oO�n������s�y5���3��쏅6�~w>}$v�盇v��55�H��f�%���'qz��Ӓ+�/Z��Hd4��O��jn=z,%��M�O7��xM���{�ti��@�*c�S���
�&�����v9_!P9���<�����O��-�(�:؀��@e�Q:S�����+�?�t�	)�B�-6d4�Ǎp#b1�k��y�����i���8����9���8�xE�yM �"���Z�V\@a��C���|De��p6���2@�����[�����b�mU��J+2.�ʼ2+h!����kN6�Lq�_�	_7�8L�7�_�-�-;�j���A\�6߁��tR���/Io�p�N�"s���t:
����{#GbhF�q�14Ѕ�_�f� G�ݖ�y�H�F�lF�Kدz�֪�H����?��ц-ᑴ�nY�/�&?N���\1fC����IE@�S�cy�*��|@�c>c�
��ӑP{D0�ڝ2k���7϶0l�q*0 @���b���'.^W�os��K�FG�
ݟ��(���Y��a~}�[ʩ��J����֯(�qՖ��2Sw�j}�.*Œ�P׸����*f)����N��>� ���y�� ��9�����m�w���3t��L�����,a�S�Ӭ��0X	�|G�/_��p�=ų�^@��WxA������`Q��3vt>,�\�\k��ր6<�-�T��]1q,@s��$���u0\�&>IS��32��>bm�`ݪs�a�a�F��2�O���KH����iQ�Z��	8p̟��#"5�\���T�kwe
���L�YP���J
����A��Ж.ߎ/{j��3���}�Ͱ��m'��[�,Ɓ���:�s/Ǆ�i�Dz��y�YHG�Gv��P���Q��7���$�,��[��g�>GR��/�z�7�(O~���瓏U��N	P�쌃Z)����H2���G+V��G�A�12gMQ7��j</��{�[�1�稏�S����z��eB��k�i��g�p/��
OJyX�l�%R$��%N��"����Qg�Jb��"Y 칂�b46��떭�4ѷ���׎� y�>\�XQAҺ'�֨(�Eӓ�����g�(��4���L�'��!{���=��T$U��Ԯ�	ӆT���p �U���1a֡�r�E���Bg�,�tA�͋�j�JArQ�����xx0}���(^Ge1nt�����4[���)��+�� �&rG��cx�h�e�#����y�u������|M�P/�7���?SX���D=� �kd�nbC�=�13P�.�9�zY�\�Gf2QCI᪡4~���J}��AJ��5�3���b3�V�׹���KA���<o�����4�W�~� %ز�4�#K"�Vh�2�_��2!�[Y����|�
7���7N[�+�V�f�v"�*����k�����y�w��؅��?�|o��d�Uܔ�����99`��GL� q�@��1���T*���#�See�a^jYZ5�}R�V����`���c���zj\����������v.�Ml�j4Dnb����'P%&��+`r���	���	�fR"��Hy�s�%���X��K��I�Ӫy�A�s.���K�GUT�G E�[����]�����^�An���"��O�>�m�=8E��2�گX�]���#�\}�)U���Un�ϖ���zj����}������G?��\5���1`�yE������N�F$�`�.�&|��p	?���a����A�!n�k�+��fYHg�����ʛ��m�k(jd(q�uӉ�hm5-A
�t�0���O���K#V��qz�U}��nߖ��`iA�Y���+�zu����Q�y�Ƹ	
[��1�@�s�8� �#�}�z�v������'W�3U�O/�ƚ��'��m.�k'�X&��P
I�������+y��>Z]��y(v��)L��*gZ��^�����}@�s#k�^ Z�����&%8��z8ā{yK�S���
�'�I�_I��a��c��g�z6��z|�=�r�ѹy�G 	�vɈ�Sձv��i��S}�1^�
tR�(V��;���!�UK	^;���D��r�?+��`�~~s7�0���LٻOT�������w�;l�I�њ��^ =`��8��Z��E��C� ����;F�T����E��+��F��iS��:�1=a�-��3'>=Q�1�,�����u��H3'e��w9-�F����ݺ��m>BW�ۜ�h+>���i��ѭ@�!f��L
�y$Ss_]�v*��F�di�2��!7F����h��.?I���?�^���&�t{=�Z]��=����&@3����)��G�b��\��qRه�sC9�R�״��a��ZkÓ�ev�&e ;���ŭ�>�y� )�4�����2�~�`��I��F���'� ��]"F/���sb�n�$R�P ���?j
�Xґ��%4�0G�+'�@=w��#���@.�s�#�ŉV+�s��}0������Rѯ&5h����B|P�ʊ�a,y�Nu�̀Us��CKCiŵg;�����}ό��9�6?�&<�ʝ�ES��*�.�8�VʁT/h���cuxe2��c�1���.g���� b����bU	����5��e��eH�y�>�w������\,K^;��:S�F��`����^Q���L�߸��a�Mz*y5���g��e4�����;�����*�$Z]���y�k��wg;�ٯ(p��3�.˲��j��Q�l^NZ�a�kX}?�⎻��v�L�|�����/@W>����s���{ti��ff��ɶ�"g0�.��ry�2*v_�{��u������7������Ϸ9�w�m��b�cR�FT�gz�J���S�z��s㼽�ó�$�٫�����\Z�r�]��C�Z6a�`���L�d�^'nY{-�cԤ_�
����R�J?�@�&���>�ܙ3fԞ�}�����̓�jӃ��#��ht��&��_����г�&�S#�~���B������T�WŤ
װI(�ZK:U��3d�ݝ�;��T�)t��@�C�QGn���NF�P%�eaW��ԴP��7���"���kioH��oCr%�x�Y��
@g��,�Ee]������{�=�sI�%��lu:��_�ĎS���e��ZWj�t��������7� )R�e�P5���+*/�״J�7>6�~"�"���dxt��E���x�[YYYM�_\+� �]�d�����<�3O��;� ���O���6!�����x�kԣ����X ���a:�����!����Zhs��!4��e�@����o�];)U�O�O�M��l��ҩs��D� )�T�/7���T����fNݨS�^�}B�=����%�彵^S"(�l�&W&��}��c5���͇�4���:j���%���	�`�g�;��kgq� ����#"p��Lv[F�)���s����i4��BK�&�}�9����uG<G��rM(��'~3'�a%��؟�}[�g�+�2��&A���$�0���䃏�����T��x����l^�w�P�LK}*�"�"]��EO+����a�pseW�\^69&���{ ɋS���j�5���OW�߫�^�'m�B�v��	~���$��w��� va�!���G�A�}8�Z��A��&���<tF$j:<K|���E]QS-�V���KH�+�sCLHͣW��I�4A�l���9fP� i��_]/K���W�p�*#����p}�s��H��+�,�)��/�:+Aop>�kd�Z�������8�}�u�,�yN�ዛ�Ү8k۱H<tbGSTb�c_��~����o��E.Q��K�î����x����A��w�-������Y�~�kUE�H�'�|��Xy�fK�Ƭ)�H0�lQ��� )����;�q���'>�GS&;�_�bx4k�e%��QGE��|��3�:ەG�R�˜��5��KUM� Q��+}�0��˗����ǅ\��糦��;q�����%ST�`��@�d��;B���I�O��b57,�鐣O�ٹҚhlP���~	Y��n�_l�XTRun;%�����&6���cY y{e��W�	ۀr�q��1=2MA~�'���Ti��\��
���8���a��b
��Q"�ϰ�76����L�.�6��&yz����3�7L��֧�"VmFw��w�EѮ9�R�Q�7��ޟ�E���3�j�P��)�(x��ЎG)K�ʢ��W,�Yվ2�����\�_o�n[>)�[�ωnL9QKA�~˥�_��L�V�,�0W��J��HO�r��t��>u{��%	+|��gG�ܳ��u�g�A�	JV�_����<���=*Xk�W����&3{R�q Jy L|�@O�i�;����i�Q�&I�Η�4�V�c!e��V���]c��+V����Xp������(j-��B�l�����n]��S@�;��/������Sv�=���?�l'��hb35
���#b�l�~�bm9�4�g'��c���t�I���#5M�Ć��ut�4�u�~�M]B�t߅�.�������GСm ���&�y�T�`\��D���W˔ ���ze4�^��*Bl�Ծ"c*�4$_�ܺ�*��'(�&��0�����KQ�����%b���Xf�r$N��0�W�C-������y���g7��+.�����<���OC}��8����Ba�+�؉wL7pM���[-*�w���5��_`YCD���۫٥җ���x=]V�]8�&vR�>�f\ n�q��@1�wY��2U�y��M���@�Zq���4 oMX�����$�v�5�pN��k�ER�
�ި8�gw��YT�-���X�m*�s}*���d��	S��h�;A?�@K���Dhu��,�sO"���ĭ�\ĝ��~D�>@:�s뫋W�@��?M�h%���'����C!�7�Ĭ��	E��^ �m7 �ي6- ���X&�u�+o�7A���������`݌���VT��&)vtwT�C\%EvzC\��k,W�H�zE�t�����<p.\ʢB�Y\�
MHZz局}#;}|Ǆy��pK�zc��0_������w�JYZ<�L�C�4��V���5&M??Bގ-�V����m������|Uyr��D�����0B�aDxL�e�r_���E�t����,C�
Z@��6H�<��I��;DwD�w<h-��ωxLJo>Y�? ��������9��᭝hd�8�}f�7ҩ�F�l%�gQä�ZO�Z��Ο�v��@�MnE�M�)��g;�B������ h-�*%!R���8�!�LEy?G�7���:	S��G3������<��:N��-��'��ϔk��̅5����ć9��}�Ws���A�/�k�l73(��e��t��UԻ�iX,��1�ji�Mj�?�����^� [G��"���x��O�b�h �R�S�	�G���Ԣ�ܞ;�(��%�'�aH)�,�d3��#S���:h�I�%�q<���������#bLl6pʑ|"d؅2,��;W�x�F���+��B��I�ڂ�@�EGw7:F�͢�/�!:=�d���D+	����R��v��9r�� �#s�ֈ��~5?��1���Jo��'rgfx�x����-#J���Q���ct}�<�䫟6�k��O]��s*����)�vt�Av5��y���r���é$|g��as���ڻ�PK{����h-E.������F�q�a�f(��y��or��_3���w�;���7\,�!U3Yյ#�*��P�]%'f�5.y/G�	��Q�ֶ�ѹc���+?�r�8�uق'���U?^}���Uɛ�M��c�� �?A?S9��AI�U���6�W��: �(�h�����s�#/ 3��OPȲ��{5�(��N�C�;T�`��aEar���홫+ Ψo��_�Y���קj8�tu�ꩀ��v�n	�����m|0ȅ9���I����XM��,HʝI�	�����B�r��/�kK����m�W�LVG^���pW�MY�y�	���v3 ���B�Ϫ>��Q���	�0�
0F�9��'��� o��p��}\�;hs���#�JH�.m/�;�0
WÇėBA͊=���U(�i��}��7�"���}z>r�W�C:g��Wu�����AX���J���bcB�����w�J/�H,ԑ��_=& ����Oj1ݪl��j�^É�7Q���kݒ�ä�b�n4�L\�����]��gSώP��1��Y;�؟č�؏C��O�`N���7����w�3��O��Ë@�Y�\񯌭���Tr�ŖEoc~�(?{dA���0�S�s��'q&��`&]�qV��
����dUʌ��䎿��x�R��4�3�"��ڴ��U�&�eM1�]E�﫞�����t���%����l��U��z.EL���bɠ���ͺG��T�C^��Ba���J�5A.Y�E�7_O�;��8(^'zi?WKEⓟjt\��6z������:�S�_s>��q	� �J$�؈��g�f���0�� #m��׊5�����V���iQ�F�X���,h�ɕ��x�4{��D|�P �p�~�"5�C�
n�u�D�H��N�����)�T��V�e,�����W!�r$'������g��͞�7����x1@�$��/%�9���6���wliP���_�d�,�R�����݃b�lZg�Ұ=���Y��� *�A�@Hbܼ�l�94v�����?l@�
���M
h������!�.|R���^��l>B�9��/���������<M�F����֋k����`�W��e���c�� R�`Y�^�U��P情f<Hb�.bG�机�o��n뽧d�v�k  S߀Ō4nl�x/.�H�*�̫W�j��x��z�¹M��tbd,��;��|WB��9����ݽ�EeU%��m�w����=.�(Ֆ
��=�ع*`Ob\6��������j)C�^G�aŷ�.�����i�ԟ&/�w������ f(��xAa7�2����
��R�3`7q��8iJN҃5��{ф��Y��@J�$��;��$M,gzCO�� �h�OЄ�V���h�Wݒ�瓀�bst	i��}�ׇ�O�a�;�~�J�f�9
��T�pɏ^�'󵋚�CǇ��7ai_K�	���:����n�m���P��J�����{���C��ZM�EQ�=4W2��*�C���V���eT��/J�6�L��%4K������~;DM��2�[���n������|�����el�u�l��ۜ�}3x����O��c��[����a;T���uД�d��SV`ZCLc�l_^�odh�"b;���]��&6?C(R�N�.K�����e�Vsp��~�Q`0u��I��0�B�����+�9�K-|+~>�LH�ʙG���	8\$*�p�TH�A&��qD�$���2��v����%U�rb��ivhD��M��8�*m[�G}ZBxZ�,�~�#\����s��Ԕ
�g^I������k�N~8j4w{��EUcn�DzҊ�@�vr#��t�~~�[����v:�����I�F_���y%���ѥ�	����>u|l�Ƣ�g���Ѕ��Lҝ���QCT��`E�v��]	3zB�vj8�^L; (�uH<:��n��h��)�!�;���(��2Q
�1+;��Y�o�}���n�-��y� ���fc�B�����(�ڱJ��͜��S�G����ѧ�F���M���G��ߗ��u���պĀ߁��[t����]xRL�D� �G�5Q�	� փ�Yo�����ub�ՍF\�̀Ӑ��@��gVn�X�paw�B���u5�0Y���=�+%�J�;��G>�aw�?4@;D�3��@z'5�f,"�m�:�ݗl�q���
���_���$�ו~[ko��-��̰��)�3�[=%K��y�����62ub�b�!b����	X�� �6kv��6�o@�hƻY�U6k��s��� �C����w.d���B�Z	Q���bwV^�b���9�����Ԩw�\w(�� �W;�E�i�գR�<���&h�GF�L��dD�����i��7����Bp�߫�%eqm��[͒»0��vw� w_߾�F����
���{�b���J@=�`���F"Iآ��כz�~v�`g��T�J���앤{��~���q,�;����u�*>��5�`n)��ͥ.x3���H�X㉄�����ܿq���V���̡�9�$f��%k���I��	����.o��Y�.�댟��1�A���W��5�8ΣI��n��c��!����½(2�G����pZ�=�J������$i�j�(Q^�=���`�e�$�U�Ig���t/��r\`��{��	�U�$�lX�.�^�#~*N�R�-�������6�*��F����L�4����p�zL �̨�+���(�r�����$�F5���М�*�Q�o��_�U��K�P^���g�&d�X�+&��ЇU�Fm��7\�j�Rwl^�ɦ6C��u���K�;d���'��I��ѹ�����5����X�Ș9�y\᱉Ͷ*�C~hsn��?.����O�����b�9�(� �W��wLE��=6c݇�^y�UgEE��-ԧ�VT�I�ƞ�FG�U�t2��$&W�/����{�Sr���.O��_D�)���[N�Q�E��� �J�{T��E1����D���U���'���\�N�1�j�O�@
���TOڙjfA=�E���+����/jC�iGza���^^�*h�@�w�JXPte�2�m��C@Oj%���ߠՉ��RX*%�j��B>Ĵ���+�B/$��||�=�������F�W��6q�M-��q߂P���%̝8aO���%1Ҡ||/������2ɼo��������oL���+#^'��lx��b���˻�� �S�oQ�f�ї��\	X��I��!�\�N��`�=$ɛw�����>L��Z�eyCY�&�$�e煜��'���ŚL:X�����w'�����L4�:ܩD�ɸ��W��mά4{^�ō��ˎ*vg�en�H����s!��M��c���W�߽�+z��P=�D��l=5]y 9s_:{��0��n�h8<o�Aص�����	�1`<�^q�ƽݧ�Hs�ۢt����h�`JK��
۔�A��/O��t�2e���(5�/2� J�-���|�_w�wB¹�k1�d�eU�%�k��K���&L��Uf�9M�uL�<OaBtd�z�A(m�J�^(C��Ϗ/��i�V �$�M��C E��Q��~��5��}�Ob;��L�r�7�p�p&'�͸�z<�L#��j���ݷ��a������
Gэ�/�*.&�঳|�Q�ߘ�����R����'
jI��B˳(M��X�
�Ȼ������t/v�eF�+��#��M�а�!��L; ��k�G&_�j�(��zE��ke��mH[��t
��סϛ��u
��]5H� K)JԘ��(k�g��R�E�!�$����]�m4�r�<a�k�շ����Q�6l���]�J���9�e؀����W�EYyp��`��q��IvS��z��ލ����R��D(݈�?��&�߱�HJ�ׯ�[�нŚ��]]7E4���H���v��&���ѿ�N4ei���-�C+�p;�_���d~���{���(��ѫ
�����׍�ղU��h�a�,��D&����"�z[$�6���T�6����/Q��?�AxrO�ܸAw#��nƨ�OǢ�sΛ��:.�Et(��ȕ�N�J�"���#r��SNdk�=`�3�J������m:���I3��l��Tl��
 H�*�r��u�\�)+b�F�����Jǩ�S��hUreX����J��,UF�i�^�w�OK�Jƶ��G��"��q�{R=���)H�~��k��PH��/�R@�&?�����ݱKbU�ؼ(�x�'��/`�0��Z9v4�� �>��O�p#Z/B�Q�d9//}�s,T�)�OGM�^	�r�T��������h�ČuM��^��ݢ�kQB�p���u�X4n��}5�t�)���!� ��p���T�����h|����Y7�$������P��/onF�2¹�x��2-2���=���U;�	t��[<�5�K-~w����Gs"T�.���-۵��Q��EA�!z#�r>͐<#K�4 u���8�~[���܌|�wG�������f�����X��E ���)g�.>h�͊4K��2q�_����#9]�Dͫ$���}�����Gl=��e-g��)S���M(R�7#Fb�?1����Gy�,�J�Hf��oa�cq���ظ�l���$?�粴��o����%��rI��o�ܗ���ߙ�����l�k�Y$���z��#8�T���c����\̂��4�k��M��0u���#t#4�ֺ����
�Gъ|�ެX$H�n�郁~4�E��~e��)�K���^���UZ�K2�|��[%�l�5����$�!ȟ6��d�F6��I�3��]K��+���x6��f2��H��[�>��L�J�Ԓo#k���<������|2fb��?R����ߦ�� �b��2��w�Xf-y"��-��cT��J��a.o�cse�t�Y�n�URZ��(:���<���Ͱ�ʾ�Hg���9C7Y��!%��E@ݎ�V =�`��Bj4��+�,��
8..N����M݇,[����b�I?�qj_���5���a��� ��JH�`Q���f�ˁ'�[V)B�. gZ@�$�HXe���d��N�l�H�����E��m����d�'�����/�щ���&������@%y���*Ć1uz�'zy�t�8i�ff9��21cu��+ճ��۫���ߥ I�Z|�[mV�8�[���U'�U흷C�o(d=�S���<��N^Ҥ��i�,�v~�
��6��@�YJ�!��^�0`_x�l��UG�/�d���i�2yeV���F��4r��������7��J��F`��4�Jkԯ��M�RP�bO� ���!�0���2ٓO��]�y���D����$.ĸ�S8����Gd]bWq����.wƛ�+2\����2��n�� �1��f�W튩�B��S���>!*ђsq)RT�B�k�#t;�楙;f�MBqT�
�}��k��k��u��.I%�vO�\�G�\�����8�d����:2̃	����co���ADϒ�o3�@����`ظ��f��Z3)�-�v���Imy�C�%�ˈ�O,��Os�* ���Y.|8�~�8�LE�ի�����c�o��B,�hн�c'uo�e/�Mt��Rz�
�N'W�g[�8���A�b�XM�L����|�R�.���*��r����s�D
 X��)�� Yn�2�<��P�FÁH�&��l�R6#c�%+�;��Rd��"NV�ld�-�����ed�i���t�>�O{���&w�?c�b�����`O�����d����TYG��Z��@W��p�oS0��t#8��݁A L�(���5�T�(�4�@�W}���w��
�ۮ�WϮ������AA��1i����	.H<��ޞ�����,�~�j���>x��O/�[� G.vu�fy3��mj�Ah;�va�^u�b����Z<an��.� 㒛������k:g7����-~����y~��)p��� ��U6x����jL)YL��~��lt��A�8��x�ӌG޽�84/?4��+�@4�