-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IzHzjm216JNeliX2ebyf9z4IRxAkARlfomphXDmf9qGdp4HvdqpbdbYYmzQP3e5iKGadEFhfjuF0
BV6NWNQ4Jn7CUS7fAH5lVlK57QhU/4MGA40pRjLbc3VHUNgDN4t92+8IgoBCLbCJanp7cYCNzu7t
mE34YnXyKRBm9PdLjddUJ1T1NOkGAVx8POSDs88Z3ubXucjA5NffKcqs/1vkv7kbks6br2Pwf195
lKuciKRzuLV1gU61TdNcaSiZdiUJVfPE7lKKfyR9bddSECSHLXtdKtd12KYgzIkbNnawdkUUnGRw
cKI6hyr2CIEMDV9DnykIINd1QKNI8u6f7g55Lg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25616)
`protect data_block
BUWL4xIPU1SAkPDbDSw2hM2CLWiG9GGgnB7SPljFkUoN7gaM/GVsHOO5TgUrB7Cd/OoreuKZ2/VU
cE95rfYw6pQwLinad6ENueL2JHLvxeNyI4qsmkAY8VaKIjQFZOPyygB1py6H62qS3uEk6DEz8fNa
2FkXroq/v55TT8Yqgl810+euJk+2LYcUy7Jn9H7lAHai9iaSDvfRTTKqRfaWA2pXkMsWlXf4Sa00
b49dgHOxz2wUHmExsfWAq/3ci1CoFvi5t8vEmjjwz5IaA5c+7MfFMBgRXds7K8UNF1Fn8xRMhNwz
arbwQ6edCbmlEEIXMFaI8TV8bCWfIuDG2fGON0hh3mZUxcfSWc5qIzl+h5BSR2LuqhGpvTB9k7R3
CTUhWHSoHEwiS4i4fIZ3mNZW1IPaEOgpi1AES0bX006Hus117pPFRtpPLYMrOH4KJvwKXTV/u4NP
ZWDo2Bg2KKPXXX7rq1Qy2oQQXYPXP6PRchEQC2uDyZpb2EM0Kz1mhDPJnp7IiR1QeUf3VXCur6R+
bwEvmur77elJDM7zQY/d85t/0vezKjO2Ye/WulSZKZl2UY1ICPnFAXSp4uDwyu+EgYYHdeu0t/Lm
k/7I4BqtokPvGguexpLLx17tvAgIZaDg2j18haidGhWM7Ftk+b4E/U4NbxCVPhMqqv4Jnh+cBS8I
5iMLnsgjOH8wleAq/la/RcLHTPVLampf74ATgIECfaFzKeFTgFGjDhpYl4FStRFEZj0knlVumKSJ
Y8EEJEVdSQEV/7q9Lv/gOl4k27K/bg9l18qvwx5I8S+xTPkQvoptIOzVFNa/IrGVwuUXLKpbAbHC
UZBfAufZuUMdMACMxO4DBJsZjgLbFsfFC7zpwE0bhQOlnOBmD/qJt/rc1TFHMHwW3Ys0PHWIYhih
qkSQDm3Rdrf8ZLPrnVAb47Cbijalnh0O6Z8NaLj08Wx/IyDA0rgCx7QiYKB/m2YSRo/iP6ZgmDn9
eCECe2ZTMd37eIXTKzJMwtr64dbjPoE4gO8P+npxVFTpXUbTAq9e1BJFEgoG3cKwstu9cV/sKV9U
eC7VF21MgqXyS7NGsxFxwWKff2A1Q37pDCFd9arSE2nDMKl+/eCqZSeX1s5lXYfWffaUBSi/ZlyS
ed5PDxKneZRmUjAT3UPWYKdQeJwyVz2UuVHb/g4YrOQznJPcUHcwtpMmvmtK7H5kjTQaf0Dl1nuV
dl7aThuQMPhwrwqRJCGK8jvS8TuGsklDHi/F1SxhaCw3cBx81xCkuh5kt+Vcx3jiRD36KyufV5v2
fMz9UTM+N4RsS3AKzmIV0z2YvAOdiJhuiy1IHq46JH7G7mc7IXgpI03+GWXF8sDS2qeSvY/mOgpT
iLm1g72SoEL3PjTXyywE+aovL72rWF90Bw7p8lZlaPALxK0RPBNTXNELYeh01CLoviCkDklvKxNx
10EBlYFOvmXEoorooPjuF8rGutcrdE5dzOTxeN9fFxpvhsqxhR/FOb509meWwuydslKg+quqR7if
H22Tlx5z0DUsWWXsN/Kghx0YqEZjkV/rAeMsAFZlBNhCdtJ4uSI3kD0U94IB9ah9K3f7gucOrFj5
NUUj0o4Br75JKe+RhUR+9qOVKN45j0ZzIaoISDphcDJwYF9jFdTBfrxZNmTS/qcF/5AhsMHh3U/V
NNewM8z2GQC79Xn98G1AncAYtMJyBEMYBGGsiJlXRK87VbsMBAf8HWGsmf6DjkE2OcQM/U0WftA9
dpJcZYIZB+ZVKnKCcJxeDxQUmMaLTHPFJQUZZkjIe7HcTxVRMtXuGRvvBGltE/2khgd3VS60K/cm
r99KdivaOhiJBXDHIKIex7gsfbV2jlzqlUa8PivF68dBqKpxN6U0G2KpOvCf5MSnbGoZ8WstYy50
KCzh0CqxtAAszX/FrCekAWeOVBKKP0MLb4oKBpU/uip0SjugmHBYU/S8iul3gPUJqGcbjkOctFxP
pOWzzYGeraV5+mp39UiE6KDr+V63VwiJ+2xox6ff+AU9N05ULacwxl/Wasls072o7R99PpDvAQTL
+3GTjjy4L5pKzIUvUjM3nHX2FpIh0c2wJq0CxhwfsxEVs7Fsdd56/xAOcPz00hIAr4lW4BHyFqBH
BvfKgiyZmTf0fkfTLpdLkAIoKl8zt8i3QRCb/z/ILc/APzjL82OJmYSbyNUKpiiZBzS2eiiVQc9n
b0WtZCVQKWtnEllW3vd5kJS13Zg4534GWrR2Zpl0+XeFzuOspOrFpAJGj4ih6DIu5LqxfqFn7WCt
H58tVOYJA2z6IZz0gJ9ehb9KNc0Dl940h/mAu6MjcWqCXrLBg4Z443FVvDlBgtf4k7+WlmDor2aF
C0HI8nf2ULNwSgxESLIRhlUesAIHEkB1CjnKcEs3xsYMjLCYJVxXG+vG4ajlu5pl2CUhs+CNT7p3
EHfpGuP9F86wFZpRBBTPimg7trQaY4v63Tk/SNiCYVKiqKGq8PVSlomKMf0HKfKDsH9HsU7WgsVY
k7l8Q8klmhY1380CmqXbZsMkmbQGF4u5yKoQqnMPvLxWfdCyWRTdXjf9oXcuIwzFsKFDT2bkV1B6
VZJuREyfCOOZYS8Qw8bG/2gb4YEC9HldIXIR+fd57b3NER33a+uZ0R5wtB5KUJRLXMrPAhUyXTvT
D9vgzDCivKT7x/2cHacXmtvITABEV13haNHF6dG9Kv8h7j5a9kkac1h7tON2FYNbAat7bX7G5org
I/smB4u3+hm+cIktYHx2AOVE2FPiHUh6e1ybXnIEGM3xyGsBSYKW2edKpCQKa5s3eR8B146TjH/c
kAadvtKaDXqdz8uCuNgPLNmUEY67OLTGNdacWQvNwoNeK7ceLQwALpg8Vz5Fgj0hj5PqzbM73hPl
LdRzK8UBXn0SRgMKIPVWwYpMKR4TIkoP0Owf3PT4gsFE2xHx5xmyRnKsBu2ZHX5ztFkt0WeQo6GB
9z+vQwcPq3pTvviNOVjALxjYO69T8Vpv5UfpBvdFHcs0xHMD1DjfyZnPuQEODx1b98wC0lsJeJjK
KgnD3je7m+7xOf8mq/1LRXOoc482Sk/hd0opWdWgKW7aJfh2HhoVEBBOSPLx6YFvytQO7WckS2mS
sI5SV6B7/3OmLB87dhBT2pUScEB+o+sbAvYc+lHV2txt8z+7CtaQY58ArtRtWbBEoQmEzRQPRZAE
OvuwBk42aILTtgr0n/26xDbwrxbP65h1kA+cPF6OwAziCt6BK1Ajf5tG0ivnFUh3EoT1JFgKR6dE
lef9/O1Twx7AR3SalKjA1mF/rDF5bIr43ASK1snPtynNjI/J9D2z/gJ3IYwvg1E+1SwrtsBFLR3t
j5cPwyEY0cMfCJy9M3RNmB0HS4kEaHZw9gI41NvAn9EsCoENKFqMq2vsCM+dh10RADTQvW+4oCOh
Ca9rq3rAE/u0+Dw9nkihg4FhJW7LSuYRzEH5Oj5D3jy2a84xi4XGr49PeOpNgSyE/JxBz3+2Io9q
YPZjL+3dRhzjdOlcrMoPOeffBmlW0KRTGSAsBtr1bWZ65ChUyNUsmuLbF1LPZhH2ovKJZDIctaYN
6fHbAq6l7a6gFc00HnarA37xTxZuVdcKcPpLHLqWxwv5R0pVt2jvVHTTAqrU/epzGDy177Yy26On
aI2zG7OyPvVcETKPZTsyMXLdCmVJGXt1PkyzBGrXts2gcXL2O8OyJNMEV2PIcJjl4H7m/mXJf/t0
YLX6UXwy/gvekvvnMSwyxEJsY9+y0YEY1+GwDQ5IJvlOAcZxfnXT1Styq3KvdJ28ToRCejqk9+V6
L6AfQnMi1j6RYOgc+RIARmrBSbENVTxia55bqSC5C3YA1eBGyUhYhScXVud/7Tf1Gekp8YhHcDoD
bSzQLVF5MSGHdVfr2fyXKM1D49CFq7fCahMGLtl6pXY0nb3F9TNbXJQz66cCLozjKs4pnAiAAbLO
f65BmcXpgXPQF1bOfw49kCbt5RbLz41z2BeNaT/xWrxzAfRnucIN2VoDDMP9BNrjk3yrEbov0lKp
0Iu/IIRqwquoSr+SZATayg9eDQH8rPWvWQcn5NanQjblrLaYoGwx7DqPb/ORtwgnVwtOslBg1c7f
l8zE7LRD3MqBpnR7RMWQe6o4mkIkKOQM+iwDMYQhEpnyRhjg3+Ma6p7O8AjpFrJsdrwga/bAVO1I
AzcqBWpjbradKxicO0r5ZEucamlRt7Cd9Idi1Kq1jJIeRTEHxkck0B4uUPgHUlhLoutGCbc7Fe+2
CtRzW5myqS0SeL4T1+s05pvHhDmwJJRWA+/SYDTKJKP4LIM2GBEmJ/E/Gv3fJNrLw3B9OCntb34Y
nKxB8tvkb2WVHDpSGMEpOBULxUa4Na0t+S8RrpkFmJ449xNFyaOj0FoRh3XA3ljkwxINrlLwuLKx
6Z+Yu1M0OsnPGwmlnHFOOLrorkW5x3qEv8XEiZ1ghzSreeBHY7Z2cCOJxWJKmYQM/uKB09dSCwM0
q4ckT++LVS4Jy6MMV7yYZad+A1e1XULEKjF6liVS9QiH84nn9YAEw46muTUpLHm0gUfFndF9yU+7
pnrVpNoOCiGoMvkyGvPfkffIpRoS7dmDu2o2Uf+2Qeu4HZAS9NSe4bcQQE/uQcdDztYjzi/0STby
85/1ykAY2qve6G886hfxZq8pW9xfUGwIZ2+wg84fXRvEjBQrWk9vOcaCzBvLLiBnvozLAWhJTHKb
2HZ7iW6OIR8m3AYb6ctFywcgKTIbsddiwO36uIxoyzWrup9t29ZpCz7vvpL8Awmf5cCfAyIu6xC6
9wqQG968p7T559695++4Xa0+YijbcV/V64TX5Po/TWSBZ72TgH/vqcGwzRwpRH1HLkVSVFDOiRAE
aDjwqeRzrcuRQ4crHfac7386lpI6P4zpvbNfH/Ab28UrEjKVk8EoTGd790KMZUYAz5WycyEN5mlT
FQgc9FJQtrWUOiIaGKxsBu0BcQD9KCfBIzJnc5J9XvHmTLoYumfObPcPmARkmR8yLdv/R8WTUi4g
cWb5fjJGnowwczj7Rkg/ZPOzmO4DC7dd4y6/A3/usV1FSSpKe4DBEIZfrdPXdz0Q7HslCAENP5Fx
CUa50SOoH2zDYh/oGMqwHjrv/ygaROHaaiRQOihVbmUmExDviGiip5iDxJJxPHC+XOFVJ2tewmtJ
KFQ6YnZRtTUBdMGMWtnHI4Qij11LBqFfjZRaHNTAE9Dwh6KX36/4UI9f48QkgPLE+3Kz0Ejkehms
xuZL/waT4uOlreNOSFZMbqn8LMNX65zIULD29mjEh0G4jQeMI5IiB4abV6UYsH1csEK2qDk8JJa2
dLy08NEkCXuGCHO8gRYuearWBQrNVFMOUEMaoA5jkaa5ED2u3fYeguddDt+A8fbbqoNI4W9AJ2DA
r5gyzlxrhCNn7MRFuUJn7u5x6uddVT77YRI8pumScuMrDHAG1bO37SnENnlm9A2en+NbaK83qxX+
uce9eYpk9BYXDMyj6har1AT+rNAXCtl+s2unM5BARlWLKemWv6hNSnjaNdIIzVCH8YoCTCXYJYjD
IC6V4lBO8+nbQwlzDu6Php9LVD6xYanqgQ6uMmjjNpVexz5tG52x8OrebxRHe5pxt0d5oN6USPN/
oaTW9FXIP+extVCWmLDC8BrvOYybasx91K2nF9Lma1/z4M42WN2e/VmA1OYAa8SZEnPPurO1BggB
OcYOUVRSWx6/iRLMPoHlVvyJl8FZ2Y+MGtdwjsoUynkyYC9tVg/5Iq2o7FWek+aFjL80DE4Toxyd
JrMSRk/HTh9UcVOBo3lspPTftTEKTBAGBcYq2z77rLqDHbrj8OS9T3ncr0usFmQ2zNSXlmOVtzda
8VBE8XHDI6nnFXDlzB4tDSaKagwU+ka9ETwrprcLbjG+TE55P0WFC9XDkrQdhXycvYnv+5bmrfGM
7DqaZ22BnOv/kfJTFTbt48f9aMw9fmNKhxhjXWAIDmFsogMs/HfiVJHvSZ2tAtI/GkqFRgy1E7bl
f3HYam3+zWVl3944ARVwiLdIlWob/21peEcO8dtd2uyokBZdYHaCMd63tKxDneoEtJ1Wqivjmjaq
kG4KL6qxJMoeotslsq0/0Y7po4v2rhMBi/009e5n1Q4KbiMqkyyNDVIrkq8Nwkx22Cs695QiDTbU
4YQVoMeVgL3/hpHqdcP2l79+BgFd0yCjMSO3YT3cQBp7hLc7BH4fawl3HUgooAxsxuU20zQ1K2DI
hn4CMabXyXRMWPFcMxqI0n0r3vgVdLVASRLqhL580bLvF/9dHEefuYhGuUcX/9xaRwryAATEoS1g
6ch+RdgH1PWcRoxW8bo6bxWiPuQoe7k74S7DLFRQx54/jHtqN29mGif09ouB0tnr0KAHr9N5UUmR
mfZvtq8ojI4Cly1novEluR3J6Mb2l5cKIomsmowsjeO5vKa3QYoqYTTCcNG0N5SaFjwTfLcSusth
9A98R55KGbR2KDbBwcY6mDhj1j1dpKcQuAE+Ex27xWq93Rh0OXDaN/FjONCMV5b6JRsTgxcOSCJ8
oKOQCg/TqtDZV4HvmRrcZMcxcJu6R7o/DACASBAdh+r1UsNyb1qA293aWl7tnaz6d5KmnmhdEELP
Z8iOczI2y5JnevuRj9yYGrsSfqrf9cgNYEWUsEkfsMVmDGRs1G2JDeFNxeH2z3zFU4xfPskOq26U
FPvUZBkmlOmc6yQmpNwgZrZHr9v/a+XfLacPLrKVZ7Y5mTt8ZQy1+lyd1xW5WX6pgoe/qCBgJ6/c
vW1iIz7yktPxl5NM3aheYLj38LwOYBXY1sCXYAMrQS8l/rDuMosRGuXeyJtPPdaSVNjlsjcZP1eV
krJ6J6YypUUlFCUvajE0QGlku6Sfs1RTy8glAIXAydqJdV3skp2hUHYW84cwLiXkoQWwREUDiMCE
pm0hOJvBHOda4jvibGN6wzEKXcz8qYjjD7AHqkXjkkpNA3MhATRDCDudJPXQ7EuSCNrrguYSStH1
ut8Zc73VTS7hmJpZk6iZh1wiCmlace45DIR/xf9wg0+lh7XlBctqt+HSFX4XbR+tXRjD9BVT7RqF
87oXxlhMjBWuu58wavxDFybWlTTNCxMiIok/bZ7c8XpP3xjDYxEi/2BsXKBiRSzP5J1L94apG9iy
KmqMqyNErkPBhjIAeBYWmwRmR9sR7axkWgzP/uxHF+7150pJ8QulHIV5O0za/o7s+KQIkrYor+IX
EzSaQM6fJpEoNwSgBryVTEFZSvU2A5hJ4LUj6X+VZauD704PqIJlrYtL1dGP6sCFAMsYp7zeso2p
8IItItIOwLctS2FBZhv5mQSvwr5jXKkBOjffaT1AgQYMApi8KEhI3DaCt3UhoXyZYjT9obst38iX
ze9mFFuJ8d1OaT6pgf0mk7x0a6plz1BD0NxDjm3D8+a2VCF8pzsv+8wxDA+qm818C1dZQ6IZErZH
pJOFeBfB+FssGLFmPLkDKfJEB8Re8xLpZXhFyiDd+ckaAtiPiQtuYNC86Eyb8tW06QuXZoYm6YgY
Gmj7VP9bib6ZntVy2L5lSH3tCwKtuN9sTiZv2orG9ZYfJgw91v/6anlRVMrq0tbeps78NVnkD0qo
bSVQoNUFcrKOSW29LmyYOO1cFDE7SwfMUqij7ix/4zK7DGvbgUjcWWhGLsArSZJFwmGkhPQjdpny
11UyppM+TCUHPRZoI/LsLaMdGYdP6qSDqpVteVPdzu+qpIYj26Aquj1VyVg+uQKIiplllRyiRt2w
t4Yqo0HmwLApgIhRRDaP5gxkIPbYzcChcooG9klnwptKw4Vf2VhixhTdPCJZYgyYdcmGAY3Oovxw
e5npJVWI8Fmk4fXG9oU2bAp8rw6tlK3G7ikYUE2PWaqCeSDt70yM9ccgVb0W46DgVYB47OKMpJnv
NSd3NDfRt8s/z3HghAxP07OHcnrL89Mqq9YBc5F+DBgjV6d+a7mhqE7yqEz449YgaMtpCVNT+NPe
uY0OhRUXuhgxFdfdhi2yztxMY8hSI135Hav9Eqnw9hL1OPfEL1nxnJi1A8315n4amWbWhzqPvqWI
4slsa/NYIdh6QFvniBHZAz/9qcLAn1NzJTrHOwiCMCgaQ6cw8Wlgb6bSbou3LPtl2FKeUvijYMIZ
iaX3Ipu33xnK+j5uigt38Es3shd/3ADztUyKs/u1/hMzgpCOEUz6dAqXbQr4nZ7K9b+JonbZAYYn
qEft1pZZCUm7Po5W7sNwZ8blV3KLAhL1rEkzDE3mQ5RSm4LZFDw/EgxSZHWNDMYpBw/zTywbE/gu
BXNCS1+YvUousbesFiPIidexw5iaxoUc/XxjckNu7r9V9JawkDfeBwsMcJ6b20aM5qrHUMg65TXE
EuxTdl9VoKkhVWqWTgwT3wtK/A3IPFQ+RUwggWvm8E0eqtSW+sXAaGjcH7LbcbrLwFyc/leYrQsO
imCvNk24mDG8d2Es6QOiITNSq7Xdl5/TJtx/VqIljopJT3FmIh4K7h3/Bxu1ZO3T/rWnpJ/DB4Fu
4hMmraSAU+2BdNbNSPUghQpQJxQ0q+iWsaUTC5pv8zY5HC9J9ZGfWrGaQ5i8deVEIhB7lxBOUiFu
Tw7MTnEQGnV7zuvJt93iYjIwJ13wrwV9uvNpKE33abvU7JAudF9aSDrhHvl/Hz2q1CL7jdW5VPU5
8pKk0M0j+Lm/pZjTc6U6naMvR/z3yTyL5ZiglgYVaZgruqmJ0Jo0TyZaxvArhAj5o5iaQT1k/qsO
q8aVHFPzjBnlp56hs03d3SLNERh4uYvx9iTB9OKj9CFKtmlxPD7cJaLeHOltCL3Byl4wnmEipf2p
gpDnVDZEVkaOTe3sg108d4qD8PrGF0E0CSni5+HPT4SNM6FCT/o39UojkAOMUAaYBXkQc7Xc0ttz
52MlZG5NjQaQ6+x8SA9SpIWNhvu5N2eXQg/adA7tGaxnMUxGVT61GptpBYWaXmfmj+2cABgHnY5h
9C0TP0vo05J6mK423oR4wdKmMLtFgQM02g7YfohO/dJQWOV61/lu+wvnZkR0CxzWoC5CNrdhp+mT
6XSrGeQ3opCDqfoTdm2DDYqliAhrtOhR+4A/hpMd4MvR4aWO62bWGdqwY9aUVV3CP4LOL5OBOo4O
ZAzHKA3u+MbabaGYTgNKRzA+PnPVjTFhiT9GtSNXbx4EW1N4Ra74FRPSmWhAENok6YGvDTvivw/v
adRtq7J2jdlM5LPVpCvJ9vkqz2mja5lIcFg6iPcoaWQezGbKhyDo0c+kt3OgUVm9RNtuQ2oaeNIn
FBDNU9TLM1Yuz6PqkSVxeu0gZy+9vo8ObYYoCUTnXcAD/5Cgjm9ANLFCHJ6/1ivIe38x9C4ggZHM
vpG/54cakTsQVDmnjlELulve7tex94++hEh7V1UuxRZA50YGGABm6oPE+t0bYpNb3SiQBKJJ0tik
ndVNzp9ohRAZtonWOTuDoXa4a3wt9TZzAd71DEMVtTVckqzHiZXx+HBiBuXgwPEieM+E7MI3+8cA
z78114+yt5NcpQVDtFpJ4Pd/OpNiLX20B3uYj+cqhob+Qr1pcWD6/1jmJBTv4/HP0QLeXVSNfN/F
xmCF4yW+lk7SxonbhbUzuNzENL7VLyWGYRfDNukBkEWSTbgMQB8WBstW/45JtzKqO3tzrK+Ojd1U
M4JWuLWbrNO/dyc9PIQWG5g4IayWfnHtEGCR0Ou/0wrCt8ubDBpfZux0JtUmcvs8Weq5YadhNmjv
AFl+rLjqlDhV4CJQsT/7gj8tlAjwtObCpfMjzAEklBj+N0ghN7zpvpSJrmB3SEh07cOZHpIpH5YX
tJKOvf9T6E3jYPNQhcQ/09Ui+HfmRJwN8roTjzCXUL9JTQ/VkLL+3fHq4wtHJl+VBlqdu4LXyJbe
O70Acplv1X10e8A1UMmgXH39eEunvURjBsDl+m2ALb+kboO0E0IjcTQum09zVJmmsJCvJKLEy7l2
98fVUEfA9xmCfw05zLsRvBlgEHsQyEqBg7Rok0f6hYPAu8c+Dffu/WDHwsWLOPO6Xi5CZduutb5Y
NMnJVPsmu2+Rmtr6R8sHqzsZZSWXZZ1VL+ZOq1usfSuHpuybeUoOVFkDZzjPjBBAJcLQa/v5brNP
rSGbK6perQwzyCQpWtF31N3CxtMxcrTL/pHrLVTKjIpTkilNypPf0Slkrs6Z67/TZqREbA/iO3+t
4IXiW2txPiPbIIUaUo2d+ih6iong6fdXp71NljTAUKS5OolHF4ozhX/wNhomrHFol0+IAS5HZ9xF
iPZOvUgQgbFKgsEt1Gp1MBZbDJPVLUiHBEIe0VSDpHuAYeOhcNZnj8HCTDFPUTE581MY5kKtTJtH
bE9rX17JeQt+VcYGokWs7K3qFKOStE5k2ygO74dlOj4pgGMXuVZjnUd6sgjr9Tn7Bdbkto0doeLd
DIlTm/MlC7KtHMmevmlgJOZE/Fyhja7QGvlTZyNxZnEPlcwyhHBlnLfuA1U3yvKbXVqSnfg+T/Te
B7wwk8mo4Tx9PxbfghMAAYV8D70Er69ijBTaXAFsEgkP0CQWHt0OzL3EZLJwp2wlOi1QogrJSOnk
kELPwqFV34xkyEI8hRYAOhAuf+zD7gvzTOvkOAaEDKUo9N77OpoSM7jtyllYCe1yo00yoqvNYXZh
k/FhfUak7iVsl0THcmc4gf18T5/ZVtjIFHmHPnAmpDYeUUTyGbEmTvOc2Wf5yL186NfP2zpV4b8d
miEFXGTWg+L128yp6Nte3bxOCuhSJlWF2ZCt+P9eBQcs5YlVkm195X9f0wdjVRVkBA/NW6BXdWqZ
UYCfU8ZoJOmI0PGGH03ZDciMdr0zG71fVOw9rzUuyI1yMJcoCecBRTsuVEzlMStaVoiDsT2lfVyO
974FvnENPODzPhmN7wSp8binnLMKH53P3zOk7/8zz9uQpuBfWZyEzVEAhmT7fy8ve2/pgL77zdt3
om69XOlfoUxwfHw4TvtUlgXSS4XOGC1nGGJsuWijJcB5SSlX4x2Us1F2dECBNikbYKupz1uc9Zjz
nF679137zRfknFL4XkuRSAweJbm7pFHtjTdSykmmeeLdD5ZUlIeSy46rkakiydi6ASyTpFtLaOxE
lK5kGe46qG7dk7eWM5DbJKqvY9+rB07I0js0J4OUHTL6P+YXnLGY1QWn2JuYQYyRC4kMCTz72oBx
Ig7J9QuiU2vHu04+RPXipuMHEIg7EmT+qYijMNkGYVv1idwLwLwo6Ok9iSuJCSvxbwuoAvRgWCE1
JxqfV5nuqmyq5lLxwJ9nfqf21W7l3gQp2tHWKhvG/REgBYxWLJObkYx728N+YA4luP36KR2Lavqj
DjBE1I6uv2DRDfsHmQ/MDtiUOY4cX5Ev6GZ3ilb4RGBTE425neMI9D+cde/xESqMHTMJQycCpRK1
pgmzfBIKEAngRV0PLjaJ3czHD6nDtK1M4soPVYHslcfvxAAPszom8yQlZXB924cUrH9enKTD2mUE
kQ57Zyw56QjfOPmRPjwBKYdLyqSetMpLExVyZdwiAv88FjJBWaKiniOhoCP0qik/OEsdPHKHZAOb
1m3FOQV3mGccIYZfmbjY0vw+5Cgza84ZHwoqzGsujIxsLKi8nqfV1b0Bwx/1eCIabUZDTjfVeDFI
1TuYBqjgp29mq0Da3a+dxsUfm07PJpuUNfZq23vHcrX21kZYXjxBClztEjeedOxHn9EaoVnh0eW2
3E26/rkcXk2PDLHvCIMBlmjPYNDitr87Y2/rI7HZ4CUMdwsc8SKSsL7uG6LoFO9ktcv2CmLuCcMT
3d88Vq1BDvrUXlKfOYGfiSLtb4p7dEQYTGQzShA/Ryn95noOd33M0m+gP5msfb3ccJUMbdHI0DFV
X2Q+8at8TmMOunuqzZFqD8QIq4+DUcuMAw0d2iE2YQ/AKeHd2dO5JFK1OEt2mz4N7BNMGsEfX4SL
w54saxM/rHMz0a62yZeQT//Q3q4CRifWSSBaBo4L0rwG55Eu9PmsdA0oNMoNhwGFkgs944lgL10P
A8ig5o2zFCHXYWr6+zgCjMSGJ7SlgWH0tj4joWWoks51+Jw5ghovF6J2cXqUJDUTkasLH3y/E64I
/IAfcWJktd2IFtgIEh+GzRq1eEWQZ2ETEkM6E6Ojaj1SAOICoQgFxXvw+pkta8diaAa0uHKCSynz
Lqw5BxS+/hUT/G6TMJq2qXh2JlFu2W7m/FlzgPHTbhsEwqity6dOrnilN2t3hfY89PphTOqA1H6e
UDJjoZcKYk8UT0NsPB1bx8ry7XUqUv0TeIXWQfgu7TqzGgtFWPRdD+O1CmLgWvQooODghqyYiHnY
2I4fSMbWMmUmh7x/aknZo8q7nnP/aNbArAJKvSbpMh4ZUyIBlt8c3w+TFg4Z5zsJpup1Zd361ia3
pH+1hh5cYHOGRieE+lulzcDCD8ytZ14dBlCOcDKt7/p1Ur66QLVrWAHAxRMOoH4NcN7YbhqNMZPs
zkjPEDCUBJjn12OWqjKsvVCs5nzIeAE10FMmdrNeHZjiVTkIqon0VEQyNseT1O1moBHiM9LclIzl
aepocHeoOXCjQydOdvcFIrz2HOCOcRrYeUMQu3giBVr+0zMhILJOVTly+jjF2IplyTtwEGQuz1H8
revc2UlAVB7wjP2SEBRhnBfREtAKuWqFki7suNoT3cM+F2IzQ9oz3lVGDnyA1Te9fC/xZsa7lsvc
lcn3x0AHJ413bFWKDp+OOfYFB6TplXqNbFNd1POXXVjiaN6biuKCKNSPg7rz9nRtW0S7fsI4kbSc
Bt7hn5SjGvnAT65e41bd45xVR0HR6+dZuNXDi0qRYEVGHaEg+Q7Y0xBdXSKOXDdY+38bNBoeiWSb
RFQx5wkqydrsQOi2kk9+/JQr7rVKD+UktmtMs2Z0kagOYb/RCChlkPQOMJaAGFqzw328lp2IMvz+
VBeEf1LWQC202UWhhJn+p1xV632ChMFLH1heypORA3crCHmUkfeWavBwEoZiKSfN9/aentEDZpib
vCUWJxPq5Jp+2OFa4HDbIAICLC45S3DKV2xEVTsFIxO8+VGQQpUzG5bCkgGkw4XRm9TmkE+ZIWH8
LevIk/kt8iOK19DJZLIgrG9eL7zkaYOadSGOdX+eAtz1TG2So6NvY2YmND24tcej39hWNOSzO/lO
+hlqGj8QLmkZzqTg4V8lavNloLeHgFB4m4+adSClVaK5JZJakJu2zIYKKpkrmqi5ENoLpnYmCv0I
Z4rKDMc5wiAQgDSEgAXxs+VT1Vz/gEt7nXZRN/YULKzRj9QA62Tzqg406QeQp/LbiUyu0ff2qUpm
RwFUOQduemh/b/IYMDYl6UF/aYVn3O52dTOh4elan5XS6qVDu6qtvgcRI3rlxfcWL54mGZTVO6X1
AKmPRNzKxRv0YBXAz0Jg1TMsAPVftvasTpAY4qlYJEFierDLZZeKWGB/mssDsbjZ3XnD3tcl1upK
X0izj58ijFHSVwUBIGH69SBnPTlX9bLTpCYq7o/81LFfT5BiZg1R50X1sGwBXfMuLCOk/JVtFM7Q
vw48hMcyMT38yAWlcPPjZXAXOVtrD47D8F8CDGQhC9fBwG1TCK6yZ3xf6A4V+JPLUH4tFBE+/qT+
U1G0TaiAJm4Cjrg7AA3n9x47RiSTRoh0lbuKkddijZlTv1/HDS93CkdjtfiScFyzeEy2opcyPkSv
mqEN4ZuuCEHZ5k047XjCY7L4eKjFEXoTZNTa112kwWV9511eWBB9qJb+VKwdiACRyXeBLKKq8mav
oru1MSWVooH13EvnTiBXLL5i1SIU2jkgIbZvHGV6YMwhM620gVGv6RnQon/fh0TOE0sWw4QR+VpK
Y8rD73wwISyaMmryJPb/vUo0fEZkawY4kXneUi4hcBGnEfZjZuQ/9jsMWKBgjFNlKXxTQaGHmikb
1YabhAi1W6d/uAQvmpnfR1n5ir1/cKzuBVtZSc+W1x9unHpax+jrQ3FkL4GruqBeGDJTXeEewVJU
LCfcWt8jbtTHw+qCHDwn/KZzYSXEHLIt541HXIPEcqBTP5OgIt/wIc03G0+rrtaMDo/EM6vQF9XT
OkmzlomCFl4Q2xebVSBwdcLUhlCoOfNHjOjN5mdUyBtvPnJ5r50DMhKOvcFIsfc1r5oUyFGRnJsB
J7bQY4ju+J32fNJvDOf347yKbnofRfyBl33UwAp0YJSEaBChBYrFw+aS93ZgYTXQRw8NCvdiRTEL
LgQ/DAnuMwsqYVQ4NQIAdvcsl6NsIc+mYQa7IbD2anKYs7uCeZdyJUm/0eHdHw8eJZdKSBo8Xik3
rHaCDpVtfF92ntMU1lgET/A7tq1ltYGGYVa/y/i8Cwsw0qbtgy9bvjF7WqI2fJBnLjHV4WqM3RQe
o6RavOEobJbmAZfpv9mtU5bgIWujKDE+p2Cqu5HJtOqF8G29EPbbiSxVNAk9sVcZujA9VtAB+2MB
qjhPUBxZ8RKYi/DFUgjNBuMqJKakjgZAKRW3bLr0bW434Okhc5dCLaNHVhI9OdQyKvE6svUSigCT
XIfKEXHqT5T8WdZM3ihE/7zLxryw4MH69veRBYlK+wRrNUhNF0IB5HKD2Ds5YIVa8o0OOpwiEzTz
VllH6L5GCRYqVa+zZttdE+ZOeOP87RxKchQ5+BHYyYgVd2j1EXHCyDMatvOW7AaEYKqvWu0b/bbw
zDroTfN29/Lc/2I5BTYEzaYY1HuUxUckplHr5SeTwh9pygpnZvgpNr51ALuJCqLSuOGIp/JJee5s
LR5+PA2Wt4u/BDW7uJs5Wy/gGnUUp6m5emfM4eH38NiT7u+3YunMJwy3Hgoh6ujeVX3bKhxz/2qt
weC5+lOxUYinDNa5oUePW6FvQxDJ0GsloXuM+EQe5hIMKpgKwMZtywu3iAmoiaY4LT4IiG9l3+dI
ILDaG9y5ufBS70Bvbw2oGdvhQ0lVBzXhRVZfqZcsQcLbsHGgvmaGD88WKaaD7MsRbZEN9uWdEeyJ
e93C6gfVCGLX2tq3Q5BF/SWAcD0MfJZ0OqoCZ7AM+/DugEQn4phhx6mFwHAPcnyebzx55uc9ZJXR
Kf4grsOkIYdvI0p1WtNSugHs62i2cXdfGCgH2Mjy8KhJlHi/FVa7gCLjbf8JOBGJul1vcMhLMEFY
OM7VwqrIodWkspGZhIpWXHpRkneF0+jN8svp1QS3sD/UgcyOAZekLOCJ3aL+bmMJYierhS6UBC6a
M+BdgrbC24A79AhPoxO5J1CBr45wYrRM32SJSk2iB8gH4Lij/jHzJP2cIv+jwm9QQOLPjWVz9aWe
XyE5Pyq4UlMGffs5iR32l0lQVbSstP0zEP29jyOjjYENZytWRU8oNIC/S5S51hU7UC3Bp3cwTl4+
KIxdOI5QsewikbwcCCTElD1JDqf0eo/TIOeL8qOfJyoxERkWL8X2oWRheCgykQ4gD1H8HBvr3dK0
vBYs0RQVLwC1UxHj11VRCdJxE+OzaTR6YhK/kAmY1BHnrsn5haG3dWrO1Y9Dvmm68mTo+8OQfH2Y
genW6p3WglqKiM6ywX/dH3nIlumdEzXBW8qbovRC7f84VfDrUnO/h5xrtmQR9dz1srzJgKuArOf9
Y63Bd7czY2FrqgRYhIdKaPiwP7YI4BLrP7wP54bqb5qj/UpyiPnpfjvFGrMM7fsQjZkmQevCQn8H
xL8ve4/tiSRT/Pulvn7OFLv7uSc8c88IdcsRqWyUc8iqfhBMe+KDn7QJ1bgvfMcfBI9oTJ2Ztbr8
OH/+tOzHSiAre9XwHiLrcJ1i24KSnEaEsUT3lhr/2JSeJsE6OwZEXn8JIqf6eDtgtsgRNFIwMWjc
LdHe8NeeUPVRZrtvXuqnXy5C8MV5txbebDHQTLFuXoSH/9EjD2u1wxRbmjZh7yg7YwSVBIx2Szs4
hQ8yw8i9LxYQn1lHIHtI10THL4dWHonQXuHQycu6tYwsY4JbH6/NgYEyferoE7ngSz206UdsXXoF
XQL6WPdWSdI9oCknUDfH/RugrIOgqAKeMZeNm20Kpr40UNwUOQJPF8tIDgQmMOc5VvSFPAQsN5J2
T12yVtrDHRTzCco1LjT9BVz9wwuOBdp7jkgGYcvBXCVNJKjLfb1wf8TpdizJyYkLcqpOoacHX3J1
zYC7uN12Eq1O8VBzgXfI4bzb1FpH+A3u+h6tl3EV/rDouCQhafBuF3nS9ZXmn+VJajlo1GYDszsD
588m4ipMY7HYyk2krrqx+W+M48rHhzvq+j6DNg/xGXWlTakGkjS5rJrF8O0+Y3lOfl7K1F+50p6Q
QYtE9XRPbGkqm2H0HbHqcf5UKHyYORlnT3y3BkVuLSAyyGG1XVV7gOOdkb1I5bh8G9KF3vU3jpJy
5MQSvcjuDMp1zF3eh6eAGGWcrIjME0Mj4RtO5aokHal6cknxrpKRNxC6kN2yEXeuC/kXQCQQNPs+
gbtDihqk3S/ePZkzRoV8qkd9+LdeU8HimjbDHRJD6kCZUvf7O8IpTl6LvizALQEW916QZazN+qMG
t0iKrswYpMntKG8pzj3qHlwoD82Qti3RjUf7ux7D3JO/zO2zIjsKBXs9hEE+F9qrySfT3my3+SfM
EE5NRCI9Jwz3FiPm8i/hsb1kTlQcEV3GijSngDGmEBl/rDMFonTsET5ogI0gGf/gZgRv1P+YclFE
u3204NnEU8ztO1oqOXQaXqNXDJKmxc2i0pCxoOY7L4yc4bqhYt8hpC0tIEDk/dJ+Hgw3jogdikuK
ua+4tLZcaLb4tYUN33FQkOtHjbUtdvxoB2Bv1DzqVedQwONyZB2xQqlUV4hF3qnXVDGxWWHEff3Z
VwzAANIfBcDFi2wj2BxPNVpqrZbt0ZYj5G5YfZLGrfqtVX4OkLhanP35lbfjZ1xWU60u7DJ/bmxY
Ka3uZ/fE5AUNNGK2xsYElY4XXwjT2/8Caql5QAWxFJMZ+IjfKYnqO+UROo0MyRA8aweU6ECmMdM2
MAjJvhA9ijvUWCysrIO8j8eYyjlsf0rFj5sbof+rrVcRxlP6BizHv7rePMuKt6myLsVNfC8CxiQD
VFh+LzS/37X7LtMLR0HdFWdgy0lt/dZtCYLKDWRPssXmp6TbdT1Uf4mp6IElGBG9n+eyIjlzF39S
JlsWMX4Svquq4MNHe7Pf2CCcHLo0LrJ+Enj/JITIu8PBwSG/u5km8c9DRanaRrxmZQ2TFaP5k6/l
SkqogD73fMMSAgAWOcbWwfuw25scuFcgzGUF5KxNIyCztXgROhbNHtFl/6TxwgCedFdzA+eWSRAM
kimHxwNCLcbE+mBEVyOpRClErqhmS7gGWUwzSMLuaoSC2LWLwx7fVqr7E9WFSjQHPuRw4fO4Tv4y
HBm3mpHqo+dwmktz3Y1jFPRx+s5jbuXmed9z745dTWS4rIk+ztFBOWF04APIjMnYz+q32RIdHcy0
bFoFWl0PKl6/iyWb4NFlW2aoNMIFMD82dwg/mop8xgubMfDO7e/ujDwZUirQiVUpmk6gj17n6HGP
g/keXhgs923IFfuYV7trg/VWsfgARAhMmEm/q3TYKeH6HVVRtHSDW33bvrU4GLJ7388JEaD1/mUV
YsR52VAGFoGiXOuj5jJg7pf/c4BHZlnZmPdfdsApYZyN3N9FdnT56kG9psRnaCBH58Fy3OPFJVaA
rjIWmRYdQk9bibRqPAoWtQt9T0jR/UzONBX40XAnJ1B/qJZbsTmLnFYuP9ZUuRcSXAD2cfV8Fye3
Py9VNathQDVNsttPJoDlbr+cUKrzD1A2h6IAjTry2B58DuAXTnqTmfYyEc34e4wVYZr8RbjLxzal
ADly+ct9bDcfMsXQw7Hck+dxhIxA/jjdJ5WRAE1aexaj3ckEp+YIJ8tDyc4vqTI+QMyilIrh6R/S
HyZ80NG+ZftDyF7L3a+b6Nc7/f4rWmd1fIPRz223gcYKeec/CQGj/lY84ga/TSmTBzGhtQSAL4wn
yy5YgamTB0GOn67KSE34WgmMq1sOPbAsxZhJJXZtL4RdRxa6IR6UbWSPfb72l30bf+8jMH9GecuF
WX2z6X9vy/3QRJ3w5caT4H2EcGTl6cpz+DzlMp8kk+t0oyGhV6pEKOk8X24WTI9uTwlCxO2hn2kF
CprNOtvIfPYeXERBF1ekoMQ99I5vQdtPaxEMjUaRTGdqRT35sBtLf9cfGA04Jb/Rk90lhxYN7x2y
41c3bUE5V0V97Zj8vTr5lHDPb5HY9ojzeRzUs2QrwuOHpQf0a7oA1mgsg/4H1VpQX+YKKwRS8l/Q
oLXQaraMU8Q7Gm1XBVP1Ouun26pTrXBoZ1hI8rtq+fZsQHeJF/IHrCRtoi50TTH8X/+Jx3ZJt9Tr
1D1djGF5YbYSrwHBLwt8fbqzAVRKddk/NmFXhTpGat0L4xKXNG36qfRqgiY7e2FjcYtYDc5u2SjB
qSKWOVlAsxwldw72vsVSB71c/5LDxUoKUoLV4Ezm7jyiENhQvY54DiL2CGyQYaTubdjsaMh0X/SV
wF/LBpUOJIPkc+zqH3x7OIw0KIqirqTzFQCgRFqlGwNbi9Y0y5JOYGnhLQ/OdwwKI8Q+YE3N9oQD
47lHpw8FJ1w1CT2pShxnpSh2JjOdv5NRFUtzLuz7i5OUgW+xYovPNOHFvG8ovglLSrOwM63SepJ+
cSoNUKItlraHEbdcyIuL9x081ROGEckUr4Ds+e2kXuN0HEEw3uuMN9JJ3Ut4molMjRkfC4Pr+qBU
EU1goBNzx7mHuVG8XWG1nO+rjteAuWbypAh9DdJx/DZmDL2oWB4m/mELvhUpnhSyX+9IJeKB7GIW
XAnVpR0+QLCff3cmdfiVtIGcVKYHU0X5QLdsyoCH1Vg2TYBYwvFlZD8fMoHvluMH+7WMrYBFGVsS
71nMin0eSjpE9vg5etL1ubROpR41U1NqncLqvidCWBW9GTRJ3YYlFn+OcEulLB5i+QHBB9C056LS
0LfzaVZaike/WkQZQkPw/FFdfkpYtGyGcNl0GL6aspz3sGm0H44y6ZZXC//A6nIqHu3OiNpwosWa
PSv5xccbtkxEzN2nu4Xfxg2g/xvw5SRDYajE0neYkifq9mtR1wtxCvPUm846LSEDv8wEC2Slpsbr
RYYj6mSy7biF472SCONpjYSNxjfRXKquAPnQWhMZ4b1E0SgPHbVppiQFpo7JwF3fb9eCy6KwUucW
WJPE3RAya8G7FySVnP/C+/NlaBaroVd1Q6q7i7TEJdN7C3S6EW4tdy14Gqpn3Cfd5H46QVhTbSio
Ty6w++rTa711AJdw9CZhftfZXZcP6HEDbLCrk46GV2dDemJyzPPynDv1wFlXki1lZaPhsSR76NAp
9lyshq14twrAIfCSGjLoSb02I5rP4alk8HANpmFrewFXzG6XFQOoe0C3uFBNfoGyrjDXUGMqUS2U
cqJjDFbREmsQstcZeQjeah/OgH2ItnVP2wxvWH9mLO+Rcx8v4+ovlDeXVefEQGICyCGigln4TmG+
wBxLU4isyjYBSfVeiwouZJ2ZRWMnGfZe47VEbnR8/JlnuRmJHrcZk4s9AxOvtczD2NoA9910mdS8
43s31m4lvHT9f2GM//SOgppfVWELbIkQVxvh4PZ0ksZuW9SNioOdaTlFUYCCMt3zjsjbt+ckaMng
XDyinZOXRCysBOfNr3ouxojRRozJwY/gpLABUd7ofQOIod4XAA75K2WeXac+gu8v8GmJpBxk5yRw
vkL4lYbyikIOQ98eNG2LBd9UakfPdGR9HHmdloi+fP/3sm2f4cMpwbkMtqE02+TJPZtcDedCT+0y
EmfklqxjAw0grutJQakLn37r19YUln21JfHlXik9h+hdjP1ICU9/uimZu5jpauJOarEBkvuxuS/C
WBREaPCmm00bikp78A/vXd+tCMAzbK+uCDgh/edMNf7Z5XdgpNeOR5FGXg9KNKCC45dk6R7SujvM
+mrPWwuaa1YjRk6AJB9BVri4nMVSXp0qwfoLaiDyXfymUP6M/yj24VGLuAxTMGy6Fha+HxDsokcI
fVCRiz8r6UeF2XqvPAG8pTXWevKIZ95fMiOurrCTYGrq9irQB2N0QVZR+L+IR8rzjxg/0bVFvca6
V8uhGR6iVaiD8e4rf+wkE45UBPETGJ3pHZn3+gmh9CL4K+9Vv0tjk/UnUg0xPz5E9MVBMMjZLh6g
whVCGxQuUnk7riWfflvlaw8bZzguad+4z6Bl29Wud6UtnyXS/gpInq0Px/d4DoJbsIh64jbEnoE3
IbCt1pz5qYhm6v72JHAJsg/YDA4av2GnhTemL87Z77Yjqo12EZ6XUlU7AXoYljevtditKhzlpNAy
Hk7K4TAX5bIxgJdjsQKDfrcvzvCr4lFVEAj/CBVDl6x3hhbSex9JnFrXzq0pBSZIxe5nfziXHc5+
+AlifnfPKhdldxfVDDGwhz6J1wkn7hGwPHtFLxG9jiz9p8M2ZFPqaOpeknLtN92sg0eXYnT2qzVS
7/pb1IpWg0brGlcZ1V5ULqwwAHUN59jI6wAcE5wxSXyzeEL83Cok0cTdkDOoTpp4Mkj9rMCxcdoZ
e5iMJTVyG4Ylulq7PWC1vogBILzff7m09jFO7i9ToFttiXhWuGon+ewWaaWIjCezwOywE3PXPERN
rqBoSqWABhoZAii3wXaRJdauzyAhsc36R4VxX3JdHmHuxX7ky1CkgmTriy4yoMbUJ8XgsIGNLAmB
PCCKHOzQItgKooBTM51SCi6SEEEemPCy0y3Sjaj02EWo0TD2KqYhYY+xLWrjKflIjt9Z/XKd1AzM
Ou1j9Sq9XVA6zk1H0tCmxaVJWmnVSLOCv1WbfW3pIj5KwEwdjKL3XZYGTDwTlREiBH8SSA0Fuv5r
WW8UUPNO/EXKda7JhK2rO0/7bo0q+t2VMy5rqJNqi3bpaBpa8gejabb4sUnrQzgNLIbESD2VzrY8
XzM5Qb7OZYZ9FngzXmrnsTnxS9TQ5vqp4ZF4ZWFyU6aOqXksIqwLK2WqVbGeI3UuXK2q3Rtm5XB2
4he4akT/7krViF56Gm6W9XqScueyCxjtkVpHZERCdmN62BVMd8gStEFXZ+0txo7EIJBmLQBjf2NH
jhhSGgpWh44xbfBlr7JLG8lAVFpfXXGvRdHYHCVBlgPyvRhkXoG8tQKh/uMPo12AexnqsED3EwjU
jI9vac3HPQg2xO4XKctUhVIM42VTBQkb/HUeQXrSjf0Hr2JkJb+Qq4r0OoGtIhq4Znttq31D6izN
WwkJzrHyBt7+H39NO6ZG1fTcyjhfT8j4vTBJ5SMHixUfEqM+1l9YGr0btEQCxCoeOmSRf+818PfX
h4EVJAj7vSgfY7piL9k1oMaK07FivobgAMelQFzjQfKehadP0zudHHsreANm+3rwL2LpYsSgUwfb
R1JlOnG8uBMDB/rTboFiK+nAQJQF+VDvf8zQ/jOk5BwYcW0DP6vwoyCMrbTUjUFInJVK1HRm4unJ
4CGCt83xZbK/YA7Gxp94F+pgXzlLbEGohMO4z6utUPriUvwKQu1o/pXoqZO1it/iFIiuPNZSYM4o
Pta0GW+y1PrvSegV6Kh82kiyCA8KcRXaDeaWRfwmPAV7ATs/pfQLMbl7IrPVnLcI/Ezl++h2pU9W
ev/DcCP+R+Hb64rGlAQIr/lFvp8ejCHVD4bXBurgCoU6DnZmc6grRs/FsPaR40AdJQNcJRDHxNZ9
xyMQ1awe552M2H6UdNQEc4JZnUSSgUN/CbFwwszW9QC0536aeiHMw2DKTb4gKnp8IlxpbAS7u10j
mLWeogtFY4xrcwIaQ1HAxir/Bg39HunmGcbQVTM+ebMu2pVytdJHMa6kFVJSH4KCpPKD1/+DACzw
WI1GHgi8Y7G21R6omzcq0t2aIZlhPoev2N8N5VYgpfLocIswFdJj0UbGJkzcmHmzEppCDd/hKuXD
SiGWCEixZ8uF6hI7JXTFG7NNUGy2RZrtmyTj2rPNir0H8KU4v5THQ90sHFhGve9AGCwxhWigoYnt
LK8KAUJA7wKyJcze4MHo6dbddOL6/CBClx55lzfNS4AAiP5ojyGe1oM8hBtrIGvS4wM2fWS+Envh
fX9wcXLXHC0VOg147lI9C5a7jIpuRIbnLZJ4u2y3kvdmWIk8H4IwQAFlb3e0aD6roWA7SxqFbtBR
G1pq5OfACID2pvEiJEN60wS+9TJO/fd/DoiuZHHYBanbWfsqdLtyMp3DmlBl7gHqzpkZJ3x6a3By
N/BLSz3Q/5Cb+GEnD0zF+TidXaWMbKQR2ToEIKqGoZeo63ZwbfuTnptjnn5aZcMfwuYyJYOPX+13
3rf3EUoGzpUWLUMcdsOfRm/Uwn/StoYPIdowY0GnNOhpqVvqEfwcP69+AjzGJavoUgig5CxHM1j+
+RAC7HakfxhDag2bxDFAehIa6o6HnIHDHCRFIJfG3jdOCYwSHR3FqnMyIQUsouWWgqPd7X7SiS+7
XsaUeSmVnH8GtE6T35Kppu7HQQygNuG9lq1CaciN1rJwa2y6u26rEruRa5q+XQVmX5/4ZJYz2WLa
AvsP/hR6ca3AJu+BycU/RLhJD0250w6a1dxNZ4CXcT48VQgDQ5KcNzdDEXGZ0uLHLHn8fTBY2YIq
rVAu6/DeMikfoe5zCgVpa+zUviuv8P6MuoMs5teparmzBvcIiW4dujKK/CT1hW3uvGiFPVINupXm
DjrMV8P5UYtE0FlmHzHJHILPKxyb8r7BynALAGJCJXW0UjqyVO60W5yRTzw03ENfnR9XLfYzw08t
l14hxCYbZMfNT+9WjFUVvzOyNwYoZAzxCR4aKIUuksbwSjDqWU7DuCh+s7eUjLSMAb5UwOkgePUo
XlMYwV0IDyG1ZhuTbK3U03dM/i3UjDRgnwUSRM8OAvxq2c8smIUrTIAhvTPEpUJACeVQ01ty6Imo
rcz2XaTvfdZR09cIsMjm7IHiAHJU8Z+rqW4fJUnuo82tgC+LaMTuYDmuEu6J2J0cbrnnEQCOvynY
F4JwgvVC3+TFCxGdlJBSB6sfMK/mOdKXg8NEmEY76a9oPryfLNLq8EV4f59wXulr7/xQi4QbsWEs
Yl7alNcXkRbzAdW4j4fACohzjO58BK3P8b7yyIAa6AU1eH23j9zT7Kn0fBVYO3Qkzr4FuYfMukct
YO9oOIEJOZFaSipjG486zebdqO35phHpmT0qCtJSnCs4doJvidtAEFDrVW9ReEpU7bEyvCsbX/Wf
qihOz2AFyXIzDnzGQ2DRcrg8EyGwP2Sb6evl2+BMo2uX2rESa1Ok9HysX19RAacP+n9zd1cobngm
xL544j6hNNw7OgyAIujFNeDW4Azd4VZQaY1P9D68hRsHEuLrhD1HtQ0nELsGDHSMj3ydq7ZeLq8m
Ck0FGzYcTU8tWfp8QtHCL2qfUDsv5bbDNwnoeRRMo9InJwXJkIjjz9+e4wcdwtnEVgfnBBuigZXi
r4Rir+EtZ61gRI5CkbukDnumrMrt76hJw9KizRGzArlbT6z7sgDl37bgl2Ok86ZCjpwrrBHAMrEl
4kK31O6LWkzfeCultTTcLjmHeivK9ja4DAkHqiRO20q3wpg4sx3d5U6E2EyGTpEbKyQZxoeBoDvL
Fed++NpgPUtHSnpC/J9xOdJyyHox6jUaoutSuCi4aTK9Pe4Hfwoo+HlkB1uvnMacotfVm/KOeBlW
mZeAV2Rb8+4lnEZQJFSvT72MLClvt2DyL4eKIvbB6UgDOCPxyhnjELTkC1cpS8WT5ZIL130L6XMH
MTWeZow3usVbBIlJFQD30vyCUZoz+mpjiZAgFYxMp860oR/k8Gx3N+1hrmerTDJWX+UjqBjfSkyE
OeUcKMHkxrQkL09CE96caRLahJgKGweRCqhMK/G6iYid9MFkZKwN/aA0ZD1SdSIPLtbo6iIFc/sl
kGoyMlZ84oSiWhiHhKVfk0jJDefKPYt3xCuYGpNoxyVQ+X5fUNSES+VkIMFrf05UQZ0A+4ubMto6
DrGRTBw1Y+fkFi2WMZIMkDUPGk4dEsKAHnibLFn+iqklu9J6Y6NlsXdm3uy/iZAIGdAdORDYko7n
hCHQzxbOOv0FCReZY/2+7VI8gT9FAnnrq9QxCCc4NvJOwSYlRhXPIMzWAm47qSuwvie+43WjEX8O
Rs+hbnJ5Ez0g0mdOxpq+9cLegIiLtruHp2hlWTw/GBvhs6dgJUbgsBKHrsoe3FvXooBWIGrsMLb7
bQK4TWzziR1b87cNwvzcc7F3JOtPeSVKa1SxYsXcdh0iX+TmXayfaRtDs4p+R3T3/fns75XaCgKX
95BLYgkiV7qBuIyVoD3X0Y0dCRmDbrEFGovrauB01qQeDYHleIcUT6TyJtoYV5+RWSnswBs3wmGf
4339gMLblJcob14lIoRdIsB/qOblGhLtObWf6pc6fS0TTxQioHvRFzy+KpWZYqf3CHgU9xI6AOrD
t3B/XOiyye/ZdlrWJqwWEQOVYuye7A8qAYIZs/dk5/Pe656qqExw9OhwxdKjYZKm1HG4YCq+OtjT
1VDZqAKxYUKqOsQdg4hjAuNpMmUF9e1ioj8ToP99P17xeYtV6ftgHI+HE0cxY6FV+IhAxkBc48k5
faLpqO0Bu2boYTRKGHEaL5uq4s+UmHLqVXgVcaCwRx8h5OtZGKUni5hpuQhdsxHfaffN9Nqu9wiz
oJZ7GPzufHMYfN0x31JheW8oS/gS78QW/ON+E7fow5q0Q0SKwuNPRaEuepth1FNkqzigHYtt+8DW
iNnpdeGQdGmT/m5EZ6xxoHcSS8kOKGcXggc9wAVKR2y88VUrg4LrSIXBAasuLFT2YYB6hA9hMzuL
PiD7ACJZ/5jDGJUI5kAmiZbFD1jkVClkv0nOj2/hCdUUFjAdYKdSYkCJbPe2xu6yk9Fv09ff/oIn
IreuzFu4fmoWc21ui1DcARVhaa7utONBKmrt109gsw+Gborc2J6NJfrwYX8GPpyvWKuwF7oTLAq9
tcW1mO6jV+BMPjfR6NJyo0x7M3fif07SB7jOtraJjVrRLO5bmt+9aUwtyaUdXDTE3SMPqGrG11A2
9Scbc+U1MBsAz7IHxvVOnLmPt3XD9CwqiF8CmoBR7zFcuL94t334c3+cEd7xk9nSaJgCX++hiDYt
vweEpTg7s6iw3K7crQVHwejNLhpgLLG2+eqc7ZPkzv2Lk6uz2omXLNvYixTcpA3lQ6SbY1FGJSui
STtPaZGngdBb1n4KbIEKKC1oRL6uT8/z77cPvus027Bi6L3AU5GTQXlvW+zcI67wEfDRGAY2hJOw
VeFaGZdYX1uc/rKF6OnH092DF2/S/v7sqestCNMd2A8HzkbGocAgORpvV1PnA9/WhvdzUtjQhh+v
a2tRR4haa47TqLAhX/5A9Hz6rpoAlpnb9ATQwpg+dj4MpMEYcDpCZrrGeK6CLOJmS0HWPoQoBTF3
HExA3rDWsAMvOkrWw9Uj249Z83FatJTuBzX21a1gzCRMPGCdmKyM80H7XpGFvu7kb3QR4ZBtOe0p
qlDQeHm8jZKOiRoBsc8i1HMSZb0VKALznz4IWuiTq9PrVHIobrV5Ce10eGQZfdeRctBGsuAYJvbs
GKP/O6G1xCNx2gAaSSx/5Wwjbd54gzabWCRsFxxCwTVZV7ChCb2FhhX6FXalJAGwUL66/juX2SD8
qHER/dJfeaag6N7Gyj2DuETf6vxg1ehsIUKDRWIT/UaM3I4km47W+j0lid5viUjl0QHUc8wcA4bm
rma2AmJEatH1sG0ZqjNItLfjAeiTIxMq5y9nABwlV65CWvaCmPYKuS6Hbi3kbdAMZ/LHc0eJcBAM
Fys4sFSKPotXfrUk8fTLT0jC3W61O9krqWNfOhkSbiJuRePHgCgqTOjXMNPXkhO8Tf3PSDQ4A7Mj
wZbkYL29RPFmmQwEFiRIrbS/P3PKuCbgLdCnQQURSwurNebH4oYc46TFE20PMQiW6LPls4X3s1pu
XiuFR5UkDZOQyR39mQRZhLbKN8Rk7VLSW0r2ICyTFfTuxSP2qVKi91WkofgR9PlEW5ywagzsj46s
cvsxzOykWTiUCU0t6te1WEoJIfeQfuXXt6EWhvmn+ama+MMPGGkBcaQmQU2uX/eF9inQqg9kMLCa
4ePTNKjjRS43DoDaqGzb7jTLriw6T+BLJRgO6tQSu7Jh6skF9vF7uF1+CuqpQ0pyL52+/qyPU01M
vIdGY3efaOJuzPvqBWOxiXVHMkMPDATOLepagNqh6Kdn8nVG3PgsTl+aHYW/v/KNk0Kyq4sHb/sR
NcQF8aspgwekmt980pleqCC0regPeWOYeSyeT8BFP6/x7X9EuPsWhexIM6KtEy4OBco25ilFhCCd
FQnOy3O/xLbW1Q+GZvrnssWx3FmAOk+GIwvOfTn/kwpwMDD1GvXYxk7F4KlzIepB7TSq8aqQ43aO
Q/rAnpcpma4myvymLG8d/KwcAaIBjUImNxHFGTCUivH2rAzcuT08Zh5uKTPErSVQRow5rVcCCdhy
AqAYF9Xfx5qNHmhtDRLB8uzpZTtbTVM3/AEs9otQLWIbdigK9lis46vpKx91RY/+XgpyHMyBG+jW
mgyEPWRtJF5EPcjij0fyixLUkfs7vPvLrKBBNJwb3wt1n5xAvfPkvTlIggtZLrTXo5Dj2uo+Ir7Y
mPKoPHun/9KfMNlQImIalqtMjTm2y47w5l6XpvrXIJ+7eJrJUuYldtYfWxtyfgHFAL3mcdrFH6Ly
8aK8jsvfePTU6rhTxNtMecmO1G5ETMhoxauQmDjRKybtabrNxOeQ44OGMjdUw25Rdgh7kOc1EFMN
vP9kJgG6MJQm07028OVGjUSh/JrIpag2ZFf0wdc9gIzqFaNS7Y6ClHOGdZ9qELvRQqxnJxA16m4V
FdFsLOcl5OHxu9/8p9TowcaPjgGGLNQJ7kXTI63DBT5HPkcH4UKuYOAwK1S53lS4r0mAGkufzday
tGfoXf1DkKYqFu/xmWmvjq626jm4RxH+5ZeU0vARC8QI5qIjl22HH/wdnmt4BD7lLs6Ra/Ptpn8g
ZpBxVZ8YRLZ6YPplmL4kVvLwBV/rEpc1FmmEOmNTsMCR0jKjgRVoBCQjGPRprXafOxjIJ9APIYCT
aE/YjnroYe0FvYQ/fw0hWjOm0dWoWaOMsK8t6UyZFeOK8Rd3a/sf2E6ejnVb5fzyhAFZpcLakst0
UUUv74RuiOHR4b+xv2YeOBko3OY1xe1V3RNdBOcoxSCQaYpaE+fPHEHMV0XdmoSyreD59jvBMoX9
erOzSsHkU3sGr1ZPuNn77+AxweBnwEvBxMjAj1usyEcn/Seih+iSC0dqKd9VarBqI85FoP8AE0u8
nt78W9Hotvk/e+MEjXkFkHlgR1AD5q7MO4WhHWwfo5pLfi34CBxFHzzj+IccDObuqR18VZWDicOT
2SeNILFDtAJTA+EDATMp1WCmmzFg9YKwPP4XBHo8P85fl9ynxG8UMPpCHd48NoF6SRnAY1DEyHe3
OInd91FXYx5FB8jNX0FUs/SDR4xntpvlfkP29hNWlvNAxcuFdKl4RLRuX4vj5hBWP3I/+d1E6oeK
dHBBR+akRNO7OYy38t3O1S/oHGV+JFPSSouVJzOUU/B8lGfQOw1bkZepX7qlITC/dMkjO3A2K9ze
ZrHvLiYjS4HedSz0cauoP7pSMzOPBanzKf1F0Buk4umlfGTrg+3vkyjKMWeiApF/OllD/WHAzBeE
9KVBJqAQzALc2JiefIe1Wu1HtbYW7KDkUBSHdJs9vR+TPdAY6T4nJBaGCrpy0C0b5OAFXPF0h8YP
1ldSmSERpvZHp8/UYmEhDFe3/f0rywYs0tyxc/zzkjx0eJGXXoJP18Ss8VkVC9J7xWsBoL+eBEWy
iIB4jR4miiSJRpSsLUO36AKNBJPYMCDXlFDjirLGs7M4HbIX/ZfgeC8ysbTtnEM1V88IUq3m8SoA
XPBO+MAZWD5yFkogj6RWejjyKBkOFsgIIV08tYD6/DVp4BXSOUaC4k9yyWhhRQlVipB2rhlNKZl+
pASeX2TY7s4Kk8WJu+dLT/u1y61r8daUGNwjATk00tg0HuelqdPzeSmvMbwEzds18PT4Bmu8hSl2
e8qtpqLifs/Xq5jWy29EpRDB/+dCi/VcH+Bp9LOz5FQIibCmhPS/FBifBNQtyaUU4lXl98+CQWME
+l0asattrRoHAQA++KrbvRiLuhXCtmmhWnMnOvSMS6VuUSDQ33mSNVPZnCvYh8rzqAhC4IfEqrWk
6cHI5qA1Lfnd977/vuPGjMQ9i/w3/nB05BgPhKD3iWCYOP4W2XQQ+PbwXcUmyJYv0IUWGHh9HC95
kIsR2oSNXBbO5nKmS1WQ9wzYloMod7zcCWnpuh/pwAsacfsW9OTK6vymAE3lv8YUc3+Ps4YIOC30
QUTMVvAXSzRMaKVhFP2LIE2A8akKNWCJge8NZ4TBqxV0sEFawuimleEEZZFZt47qF/rJ7XIg7upB
i2TMtH+9aN45WBxFVFZYarI58yQvhV8Dp8g61xSQrUPRB0RvQHgraZR1h0hgxsrf+YI/rkz4JPhd
8CrQTmY89epSnFBHngbzHviW/ckaI2WMTofQ8yaeDoeqXI7krdT5O1fTS55OJfzLKHLtqkRQBhT2
tnJvIevROCvLZBbpdDD9cvsIaQwu8VUsmNJ10o5mwPez14EcKV2+W8SdzGxkVmefCLNegkNOfF6G
sRHhfUCjOFnTIpdAUF07sjQK6JMgz61nkmtSrmrHFwA82BGhDaZuQ1byM64Fxkg5fUKBQJrRxpaK
Swte8kgF4GjvCID8606cf8ZRe47V+oRlovywKKZj3s5sqOMUlZM9u16WxKLa4dPYNy11aa/CriAA
U8NFKECNZm/vD2NIVWAMeV8VBbyRW2UwljjiS9QLkzC+NFh3eAF6H7QssVkIrTTWSX2FFtIXXLq0
juT34kZd/CIckth2G25J0zVptbUphXK2Xaqn3XheZtb/E5uouRUsjftpVZESfnrXXR+CSYVZP3kW
Nov6XwxgoIn3VZjExdb/F18/mDcoS0HEjf/V1MTI52J816yO8GJO9R7ERZ7r9qcQv2+OG3uIfblm
j5wLdeBIXDUME5j9QWLpdlFHtrpJowholnpzjQ4dq9+ZyiCLYXmV+GazcU8q0rurn8vg9VVCmRDr
pUR9ES2Vx93EKgknMTvh2srX4z8+bPdXHc0ZO49nTR22J4tVeVxCXgpsfjnjtM+lz/jBNfI0lTKP
uikEeLwahuYaNhSbSDGoBT8XbEdsVj+yzA2GKs38XEArchxZRPz4pQIzOGedWBnTbwW3nowxqUf0
lrvdJqdjnI44FlVJsmImig9lbjoiGXc5L/I/Nn0cBzUnJt1MMszF9TEkm2ApYwblDGPe19t5J4EM
PuLltDrYUZ2IRzx7jk+Y4NJqgSAIZK4NwbxXOb6GrYYG9HP27bkZy/OZD4lS/mmnTx4a5VoPI8fE
QKQL7LQVaU4ttSd5pDLPGxTB11aQwfTAz3rFhO/MvyL3jxsyE5sKHwrVlOlhX2o5Hk+L8vE+jaAR
+NdAakoVQglAjx8QpCUdYRuZZ0dL8hOz+qGBejnGLfwSEaTIeG6aktEhy+X7V5sRHRWLrMnmEydx
yJTZ1Jmgs+c7RHHTJ4PUrMoFIJtj4amwRuZv18Gp+IUs7iVEndFsCwlIUrT4CRPoHiws8O6ngG1p
YHZcSd6n1s6nHAu7MfGm+Xp9yNoq6wphfo/ITh34RZmI48j+lbC7hQ6xT8bGHFKHl6GOwGiXrmbH
xmQDJB0hPSkL0evTxuRrf67OwdJVvrpDt7TTxLObFJthr2Bn6JGeqZ0Qkmm9CdI7fZeee26VbpAe
qYSdqpO0TcYyGdvbznBo2Z5ISXuBi822uyCBoPTUsfGcSaxeMTuU1RNF0s7KE4qZ16M8D6FC3k03
5YHYoyAtYMGXUKejIQlFkGawqA88ayO2p3LSw3OjUD1yNukQyuAz6rQab0EewK4/FcLfrrSZmyzA
yx9co+9NWqI3FuCtpbo51ya/sbC6UmSh4St6CCusYzTHADqiRl01Nzisik9AqoAC05Mz1BZQG3q8
oFvOamAg+6mwqvEutECfuLKxJyJXrOTScf5bcQsjUSIg7qV9Rx++KOyu9ZzCFUd2m0lrhgiRwNnR
b/xgGcRl5QInOMOzh5dSBVIYi/nW6E4Px8894BHdObU2ddPBghm2sp1oBrqK48wDADix/dWKU7hG
LypW7u+hJAErJzx9nFfHPOabRNpd1MxAyViI7+HNLWKJn8Z/7Dk6ZfoaSl4RLiqUVIEReEMVGwq1
crl+jdNXbEHvhHeOmZAdGVcFRhuAXlo0hhkPoG+I9VqRMcf05vWyn9tPh67yFmyfx7SnoCJIhMpy
OomW0ytSExYcx+9VpvMzzBkJJNF4FZEf15dX1cO5vqbPm9OXdgUyOZ6AzBsYQJezbmvv1IhJj8O8
Gnn2FYOXd5xvSeRwrD+TVvUCkkKJ3nvo7sMc5T1m1/KSE64RJKZwMioO5tzWRiYoawOffq7auUZU
YH9NCtkFCNDSTP660wqKlE4nnfs3MT8ZQxRS2sXm1IQ0KFntljRG3HwIvh99DqrE89+9GN06wu4R
O88FuAO9GJo0QYtmax9hScrSyaCkKdBmiccYJJimltNqBVDB3yiLwGagyd7PmG6utms44wOy0QaL
8PD5RHNhnO2VIICVfABJw0oWpjgNTZ5ok3CELQWReVxNSXFWAtVh7nOeophXMQGzrPmMZP7VycwE
U9PXMl1zdCknxFCsyKk2qexm+g55YpOm8nox5tQ6ftd5ypnwWNy5cMgE9sL9fSxBeEAPNrgVoKQY
qaJqdjbpnnqjFfcDYPWg/YL2bgujTs4D5O5P52OShnvT0CpbPIOrnQxhdv0LdlHQALqkoGvsBKgp
3IJGpMFUsd6pf0Uq/e544oNr7TCutByPuIPmEi4lELeE9M7sUdn5U94QeJaMhcFS5VKqQXS9F9nT
wOXSvpOQTWE14PaJuaeV5Njo1PG7XzUKfrp/vQzDjrNBxZuP86Ak+cMiAeGRKih8g1gmxJTmTdr0
G8iQwqUwcCkpjXlcQnJbhbP1KBXiSQ+QGfLbRPrXqxQDJtP89UlJwa1Imu0fIiRQ++anzDEp5Sd3
/ZxbP8PASdUiae2G+c17h8MucJxIXep/oXkUdomJBx4Rdq78QzL9hW6MJ4jjPr+E3SJlWvCGYqMz
8jhR55Aqv7EErxheHx5d29112lDPtDJXMpIWt/BHDNbYowFfpf5vbB3IgKFxr/MW55bFWkgVP0uJ
k94rmooZ+N8dCKFHw5Ziq+DHiiLuKpBghR5vnz0qYL08WPd7XdL3WJQvbH6ZUJwtbOcCyiXyfbcR
2db6e62zGxfhAsDZVaxWyeeomarUThInYiJwBJrGv+5y3VQhWT1jRAc8CgH5X5bgXZW9LetDYbp1
5YYeawI8ZB69s96AHxI/5h91BoktNCDSBeILMA7nAx5xfHjBd5x7mr0Gx+KMt+agXf6Gw/WbtdW6
sT41h+J7CRqj6sLdqpiYssjZOkKph7UWIA88DVNYD9qhadLNd8ApHG2bvLExzu7VuNLRZl4ODWmV
Lm7gav6MQYxlRRY8fmXfWTaOmUD51ubzxbMn8pN5F833HcoiH75M5bGzkVaoSdHQfMuujdmDu2e/
0nkENFva3M1jU1wU4OWbPXScYk4J1cvbMndUtFFdjLDUpB4RUuHAsv7m3AV7mrYsgGfylHfBTXuN
PyafurTBR4e8zjHuYwpNQyd3dZZ8cgerYg8rgRXt/wDNwE4KJqs/SjsU0yTodvRrno5zI545vbxJ
tKpN+FJtqNhsA/4QNw5WUz35TE7ywKlJh9Zyzus+5md/shklZGJMpcMeZhOp9z/Udytl1TU1JEAz
pZBlryhlODO6+YbNF7kuqYBLOqsND8KN+lBGqkKUFxQ0MHhYPINPYoFxJBmk1K5GD7ZyseM2HXcK
5IlO9jHIAnXfOanbrCd6mvI12IFPMBiO+UhCZBFCy+XcX8e/4cgExAOzjbZkzfcUnrUmrVogyuCm
Ag2J5ASr82E0W0+ZCvZP+Xrv0QufJKLYAJdpvdIm4DAmu3W26hhSMQvwLFhe+i8Sy8h6tLnvZHhy
edKhMkojbHP8gNdcIBO5QlMFBLTBS5XuovNQjw60EX3usf8ibS9pdBA81n5SnL7xnHSbp/cU1xjd
urNjhnuEZ6gndtViE5lpqygHWK1D6DxaXkfPrgHNl2SkU+s6Hs5r7zgJM7A4KW+M3S/9Bcq4tzKy
COfvggPSu+aPUWzJVIsZymVsYGmvomVV+iLDgr6MxNOXdJCTRcEeoyL+HU6lJpLuz9OYAprZGvbk
Uaxd3yC5thmX1kwFDwe+2Ue0ZOhqS4YkqdrQqD2WAnh07mhkOPSoe9ydAVihim+tsK5c2S6TCAyN
djKg/5WlLzsyWDoXl2Tca/VhMvF1oVWGIgx0fpVtP1lcpQfampHHpWT62jinSKreegaI3B5jLCY9
T5E50dKft+PtGRrDA0SEFqV6Rm+LpjBIvJJD4P7+2blUY/bA2DzvH26pRNHEPX4z7PuDSEcn0qhe
7Ot0AwpVpOyXUYHbn2QHTIal+erjZ+m1kPoruscnX/1iz2iELT91gIFSkfKtq8T1JSjFNz0OFCMe
hh5IyhHlztUfjOEOuKo7cDjtiSij06+QGbyQA7sK1Im3AqXFVwR1SKzneedp0BiORFCBO9Iv709T
7zJj4t52rQtHAi9gC5KHcRd6psHZrLP6+fRpykQMyj+C3bOKebusqLkS7dxEj89JcFjLQy/2XYr8
m5q2G5Hi6eWhhHV3JIB3AbxtUr4vzdXHneyaXktde/N6eQB8VYzmqqagTGuVf+hSRpflpjW6/pNN
A1rT1YbwkNLLn0XKOOj5m9QC/uGa2eXBnkpFGnWSv/Z+SUwQv1e3NSNpiKdfDBSbHZXVPGLrvtlD
OC2GIjd5wpXXTNDeEGNaObDvUpqlG7URaHxYCxA1t4ak59p18zszGRrBV4YNKz1cYlHVAFFt44iu
eg6/ut1snNG1oxwcwWsuD4owo3QmummzSlnmLekekj9pACDSBYexegGQHoMLsQgQ1VSrWZop9D7c
VxoxQEJ4s0bFg+jJ2HfAVFvjbrMjPmfn922sQR0UzHU0fDkbK+0gAGcEXBGpFLLjLqFCbWMKUoJ0
FUU//OM+1kKcujTkrn6ntRARz6Un9+Fp+C3bPxdvRiNSw8md9mGtiU/dO8jJoi8fIFaH1REFluoU
tRSJmbZl7OFKc10RNswtoSG37P62ZUqpHvhZsMuQUHwfNmgrwfL3LGhAIq/WimD+KTx2AUXQR3Gb
SxuvNZMdcq2+f2vUVTSCv8Z9ueHw2RSJxIwec3Gyml3vZ7uQKxbBbNjPQqdrRWTl4dMh/tp5XNor
bN1i/PIofVc+xie9Dvay31bK760x8d5c6xN1LX56/+KRPoxcKEl/jGIfgpE9CTmba8+Z2i1yFpso
OFa+DMIVB7Dh4OsoWButjXQlbKiMEpYwfeEds1lYX0LS3fxpQum5a9IDfELcxsHUgn+bWPjGwm3n
GQHjgYOh/rkLEIyfnWWFMLo14AVitl8+51kbZIU0SQ0jwZaHlyqpuauCswmLJkPCemTAValstpza
HQ4YWhfhyI4V32K2fNNNIEi3Fw8oPvDTIUU7+YjcbMh6SJP5mpjH9vrF9gm3BVdqPIRF5uhq2TMU
4EA2X1TJSc8V6woujfpoq5f0mox1KuihxoOX9XcgOe3i5YN2OOec7OBfR8+y+fNGbXxnD7jGPlDF
PHlUmxjph5HXgmn0xtXY4mpb5Vr9nPaGceis4a7yliSgu4W2emTHPktRukTntjsii/GKlC+MTjhf
v2a3FP52wqghGZvD83YgY8Hrwa/Ihe9I6Mus86np9VW2zGXNrKAAWPckTM9/6yG9SazyYeuMcgpa
yLSyeEaeA98NWvhMkdqr8niw8jnNgp76LXrjcm4PzTGJ7rSOSkySe/w7wGmKefJKpeyCrxi+m783
PGqrinzVuHVjNytlWjYzIs3cizkcrSZXzUBOgRAW/BqDcdWnleQhxJzUOIn0wuH6DszfCHWejPzA
a3kd8WhCzp6I/FS/ryCgrTF5cTYWxhZfgKYQ1hauTpZFxs7lwXlV7XxdOrlHao+ecpfX3KlmR3gH
gp91Y8KhdU9M4MYWlk6/HEfYCKJTaRE=
`protect end_protected
