��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?����K����|q8&�1��RG�|
������p] `'q�&[5�#̣Q��jE�������'+���?&�������������FN��6���� ��u�,���/�օ�q=S��cȅ��eI�pe��0�/�0��-�x��D+mgB�<���̗Ȟ�9���8Zw�X���H8���DPc̆Yu�c���J��a����f�^.���?�"���IiH��x!��q�`�������R�˚��J��9Pb���ˈOR��9�n���<��O��j-��������W �0`	���5��ep�1	;,�[��]���"�M�B��K�ۄ�Z���MVf.��{�����^Z<��7���WZFæ(�W�:�hEjn�Ė�^����q�֪G��S/;�U����
��	�S��Q��bn阽���% q�32���"o���M��܋x�e|fa���S!����[l���F_�&s4����g'�6�|�'��Ug��#3}2?0��ƥ�+!(g�y�B��"?�j�_?�q�o�P,�x���RH�U#J��z4��ԯU ՛���!�>�;~���f��B���Cn�-`#ƏQ�'NoT�Dn$ ��T���M��A2�`�
�,�E-�T|�[���؞!���:�bT�NU�:}�&+��v�6�7��׾l���2��gu?2����z2'?�X�?���XW��D���H�|�g��W+Gyn��;թ�G87S����t�_E��E�b��%��LpM[�=��H��Vy��b`ZB����� �QS%�w����#�q�t����yB5�X�'&� h� �VbnJ�O*���x K�5�Ni"/�3=.���˷��и�H���PϻфO�d�f.޼r��~����Ǝ+�k %�ik�;J9�fֻ�����,nE؉�1N ��␢b�lPZ1�
�K�"�)l^sU0�u�����������k�[��J�:�m�~"H�jt 
�Z=��sQPYT�S�<+O�!�f�!�rVRP�IO{A�j������u{�8�y��z�n�2�4��>2�(�/�ы<\�_c}�O㟬N��3��4l�g��|B�~c��}6x��&\�E�>RQ��Jcp(�������;�H�j�P����	�D�F�-E�n[����#�ƹ\�0kY��M3Nf��Z����x��[]����f	�'I,pX� ���IS���/1Qd�6����%�t[h�����>C�kLЗ�V�6�b���:�cϻ�r�2�t/i̮�ҜÆ�����{֐٥�C��[��Y��X����I����KEH4	���9qY	I��]��1���~ˑ�4|A�l��Z�F��C�2�e�!���ฐ�d|P��V1��.шN�/���Y���-�,�/J�qw��Q�ll�I��8Rέ�f�BK� 澒X�Lۦ�����gS��d���Գ���84�*`ǡ�2�!����0�Z	��N���0��y�w�ip�/��L���mv��	��bO���B���_p\�}����.�������AP%8���ړ�e(f�^'���i<��������}��rg����'nvw%�������$����p��V^�TN?�}��%�j��y���%�E�v�@�{DF���t<��%/�|�2ņPm�s*8��v8��W�zd��=��U�*�"1?�����!7�T�4K��7�U���ba����0T���Ո�ޠhm2�N1��\��\C]Pf�ZM�6��C3��#/��~�X����V�gem�tt��I�Ye�R�u����:�8w�!��C����<�	���0jX��Q-��D���1�#v���D>��U�0��y�q�DI�z_�$.d�0���t�N�,��0��>i�a��V�ݫ�#*Rt�^���j;]5K�2����k�_~�ք��y!����*l���2����ĵ�X�ן�W��>@��]g�˵ܹ=}�Q����b݊�^yL:<ؖcS� �c�ς��1� �O��}�zc������`������uW���iݟ�<�a.(��ww���҈�,o�ᳬR��G%oM��8cm�{�S�l��ƴ]��z���/��}��$�h�TR4c9�F��A�]j���2��8��	Hq�P3�eC�U+�F���j�\3��S��x�0��b4wGg�<]:���VW|?�J9�wo0�K��a'n@ע��́T��,����8�}��?{� MDzFW����}W����w%+ik���,�~��&��r8�B����mG�����_��
��ʦg�}�[�^�h�����������gA6�v"��>"��'E��Z��l�o���7{�hτ�g���{��"?X�b�ǿ�J�;F���A�f�JaA��^�N��:���qڏBG,���}:򐴸�X9�kd����d�Y�֪����FXo�� z��_�P�#:�r�d�
�n<}249�!�J�������j����0�Ű
*z�D�	�Q!h"�,秆���爹���R�8����:Y)j|Y:��7�Ӓw���e�!��h�_��m�Br�7#��}�N)��d5������g��Z�#p��l�h���n�@�3j�[x�ZuGiC����x�!;k��<.H�u����c���wa��LPC��/Ҵ�1O���l� �)�����7��<dԾ���N��>��PJ�񩗛��a\�3ו|�N�u¨����n����{�7jY��x�
�����-�UB����/J�m�x�K�ĸ�4I��y�����8}�}�R���^��&4z�h�?e�zɜ�K������[�yA|D �e����q���r�2%��W2�IE���Id�h��t�#8�w�*�Z�S�̹�ϐތ2�`I&U}��n��O�T��h|F7����G>����ԛ\�(�3
8 �~s���9���G�D��wK���z�J���M����nϻ��M[�O|M�<��ه�#��G�"	,���d�u�Ӷf�o�G� I�"�E/����eI�6�.Z�l�eͳ��Y�$��$�~�Ho��윻`���!g�,ocH�L4���;Pf��2�t��[��t�K�v���W�2:�jx��
� X�zW�M�3�.����R�:沭g��n�Di����Kdj�Dq[N5s��w�lНt#01n�BǛ�8n���R��v�?�φ_�("����tҷ���'hg2Т��~���9v񒰏J��P�mŜ��o�g�DrKzfq�' �:jCM��S^u��%�;�a�؄R�,S��j󧊝��c��H��@D:��>ՆY(�������{Z�:8'v��rV:wP=C^����a�:�?Z8ϴ�پw��2Σ���,�.ܥJ� ��=B��j�� ��a�=�h���3��	(��,ЧX˭Qאv�7C�%�Y�O��($(,����9�Lw�*��t��ԩ$i�	���%�q��6&͢?˾c��lB���Z97,�ΐ���^-��5<�P�3�J�*i�1���#��ۛ�`��H봶H7�T)fy-&�6�g5�⎘<ݴ��-w����H����XL��89�c^(\�aX��l��C�Q��$�d�ᧃ�[�]-g�d�f�a��z��o��-����1���S�5�1�W�^[����peO�)}����>�3S��=[]'B<�8���@�m����+�I���JT�6(�b�;��k�o�hܵ��K=�O�jw+�~�єZӘ�%񮷀QW.��&5���< �k���0(���ê�z��>&��Z�f5<�Vdb����v�5�&(��Ko�Q��쫽2������H����oA8���E.Qͼ���;��
�ꦓ*b�^v��IG�܆�7�K1V�l�K�F�:�|�n��M�w(֑B`J���d�J����_I�R���A-�AQ,���@*$#�-�Eߎ�deR��X�Б]b)ЍX(�C���T���1�%e��<qu~�VW����XV�h������K�����Je{a-ү�?*Q�;��D���!ݭQ�̔�g����;��ލ�nD�t��|���Z��m�_�3�NսH{1�� Iaq�Ϗ&��.�C*�����b�>������1v���~l�#��U��Q�.����@���i�j���֟2��{�I�S�f	���K�b��? *�T	�/�^F`d���	|
$��[>��g�臂X|�~1&�̠!a��W�C�φì�