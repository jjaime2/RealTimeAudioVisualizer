-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IHBy/zqNOwfqfbNbCqp65DmsKkCUX22mX9d7Z6qg/m7V9QzJoa5m6Cf8JtXBgFM/R15ZAk/ZPqUQ
AyFJZZfzA+ioEPtzZHrq2f4VauMwm8iFQPTXQ4Ovh/t6CIjTGK26IpxzvlziL+Le9Qa5BjOO9zTp
zYkDiJe6AXwcI3/1ILO64NggKXOIlrZI8vHvoG5sujQRuly0W42X/UoLA7g3pRjREf6JIKStGtBV
W9UpzkrnUMEI0/HbuITzIMrZkbBWAd7xXTV26+rPZXj8ljQspuoqguaYsHwMbzj6McNkGJEyAAkS
fKhc5gaeT8sSDd+wS9UkCQonY5+6kvBQYrleqg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11872)
`protect data_block
d02q9VSYu+LBl6kSUTGid5o2pgocpvjgUK+MSpGitxHq1ChvaRC5mehqqgBZm0fmWt7abcPe/wyS
dKrQ1H+CHIAwA7ZXmRA7x/wMNX3Bv6FMPhLBYb/MyUoknf8yMdAkTyLJsDaRT8uZZ9FIr+WxTPy+
viOKdXxQdMCkCRjcddDHyNbmGiIQ/k4ONkJPspqT1ZUG70vfJKLmH0qVRrjeHrEof7rjTsOnCx8I
6ONa9m3tq41H4suA3+KUfsO1B/Ol3STlV2sCuuasjJeR/A1tNNwZKzsp2j91h9v0bRfdSPZwEOKL
lj2owQKenTjDmg7TfWV5ZFI8UkF0LGXLNF1XQCJzdIkjWmjaKY7U3cnz3dYcFwUaK5AJF0mp9OHu
YqSFrni3av+Evaf3n5XPfKwA+hjfdslEDNM1VfrDQrecJnEF9XsXDSbMei8PnQJv5CgjE1YwLxSx
2KvpQ1WOvaPVAM6hWxbcTOId27EcAW6PtBFBCW8o6BCdyMNAWyt4jobqkuMcgmNwzlWrKBrmOpAv
HfqlxJeCbN7EMcUKIfIPg0oNJ3eoDySLzp9+GkegS8AdzcbIAXDlvaCARpEvrREu815pAiXIaTbc
TZu92sI2fRMyH6AzXcavHiHjN3yutoVkrC5sNF/EGuje91FxOKSpf/28++UWVczFlR6/vC/0P0q9
Q8NZVkK0hJ571yGBu2FCUFgzCd9KtywVNjSOtJw/GPCEbz12HTEiC+N26S3uqlBkDGxmVovycl+z
ZmOIjMSxRzP+Irf/QjKRKHkFgK88tdtSm+e7hrgOU02qgelCwVvOcEiIND3alKSguLsKbbnX+yfx
k2yd3EsBA5nNnS9cI2Y6lGOcjim688iqcJeU0Qk+sSmTTTFmD27QDdZtCxH8vWYgeLrsjZTkw7zh
Fo56FmJguHqSi7dO+EJV71bqDITw/Rr0unvQL9rRe2PCJ2v8WEv69s+tSDNgTFb+4+nZ5y6FM4UY
vsdwrY/hbu//5UGx6dfOWQQMetaMxiNX+Jp4/GCFEoEovvMfdS5OmBGM0Jl/9Y6xyuK0MM0FJ1QZ
I10D6KR8oKMkU+c9/dwytF4B3iAuuWa6x0Ak4UEB/8wG2b5SQqcacqBbPJ7VTf3krhbimTR50NxU
GxrD138qhwIoG73sO64KpKmwmfXazWKbDRr0Oyaho4rqBOTI3cSApZ2TlI9i5pv+t7mc3ZWEVe2f
HwVeLm63Ce9ULnJfh4W77gc0s52CeT6jqEmvxl/z3MbMOwxZITD+h5rJuM2ST0VEpIy8oBWNSQ81
l9eYv2VKwcD+i4j9ilzCMSvy/iaMevKNabRBDZ33Pp8ueSp4J4KsRfFUU0fPMhzM3GqyeUsSLqpv
S4YYtkwHNYrCYpcqzPXFkZaLt5ELiJldaxfGx6cyIXdRpL2nCCagn1O0zYdjeM83ebVlpAJocow5
TnDq5xvYknHgJGzVnDN2L9RQfrh5Nkx1Nv7QlEWRtqEr0YPw++bxgGgTOkiZcQy20qCF1ItXvEqB
+GTVZlqR2m9ACV+hByMH+Ahduatubna5pcdOKo875OhMwMYEIiYDeqgJ3FlqbbNh211HQ7Dm5SZH
G+z2/OxNP4npRoEfiMGOUpiZFuqzgEAJT6dsN4Aa0tMx8ioHld3Kmp/mAo8OlTIK5/czZCYfxJwm
ZGykND8e4ygHroz5BCX/rW2RFLR7ChvA/kMR1t7bsR5Cm+WLZKNsqZiwFNtfTYIyoiJB458n0+S6
/uxRH06VdAajVGNJEXJ9OBybS/i4sc3pbrMeGjqqrqtcDUyYate5QmvfiXaktXrMAbntrd3+rFaf
EypwQErnFAouBhTXm3Je0ELROcMzuGehe8PqmyjnkKVJL8U2DZlnp6Qv3fcl6Z83yBJh11vl3xCs
4M0AAbaWrMb37oH9H/AGj8ecCdz4sZ/tScKwv5v7ObKJgTXNM/SY40/XWPQHK/Cn0opAOxi8u65t
5td5U+m4TIuPhUWXG9BSBttQq/H3gNmFGe9kh1CiQTzrEqwpk5NZWJkuwSwOhT/aBqIIObA7jTPu
j7awQYOUBqKoZ2/ef7fKet+iDrkZ8kjY7NCrwvhvIy5I5u3wmhkokdnvPSLsqM20UqAxro6ucWF5
mUfH1uO5Mcp83g+k4HNCtUupFB+K1MVyW61MZtCcwe97PNca7IRb9uzTItyPOi4F7jHSRciPnPV5
4TfpB+8lK9EujKENeKGOnAWzrelnOS2C58hR60+9pHwwNzMIiPsYwCppwH5Egubj89RFDzRDw9FO
AVEUA/oN7CJP+UoIHimx91KavnmG8MetQnFeYHlUc8wucDSWZeFruK2QA2ZH/rKRZqRQ7+sqw8jT
efJn5RQ7nBLjotqfe5xKS/KJQPuw82CrVBwmUJFpIku9Hr4srAi+g4zA6Rla6T4mhn6ST5lVAGi1
oxejfTZHBhOrc1dqrXTOF9VkGtwNtApjjoVZRL6O7gqkit2qk6vv+w92ZssgR77Jbs5dg8JOfjuP
9O9W+GUScLCapjHHsKdGO1d69YsCavtSmv2ugthijkz8sCIo7gTkP0by5zzl/O1t8UooftSl5zkz
JT6nq3syCU/Y8bxPcMmDO59Cidy9dDKpLo70PKhFsADHLUDMs7YkGBr+PVtUuv5YXsHz753JLhJx
rn0drgbx7eUeZx/MSOL3EnC3nljgtiW1fAYo97pwtOSh/KsllAbRgavyu7D2c/tIUesbkHMficTj
OhLcz+2uBVMZyJhQULRFpfXhmqv4FcHf6crIpzR/z40nvAQoiku+yYAoa6iCgkpjx19H9EEkFNKb
ojypPqg2fooAlIomeGuPNnRSpslcrgF7CIeLfmdPBq05QP1AFBd0I6DGR4FD+TLUX4Ofnd2H9UUW
HYKJauP2QREaD9QHFJbtQk34BvuL1yBMkrrScbyVt2jAdA9xKmPo5Xm+Ke+Xu00Dg7ZAC3Da3ftr
5YuU0gnvx/MnLhME29yQsoeGBXAYe/n6Z8rviL7+sLhMYcFbiKDYJ2tg1lK5DcQGDudLALvlNSax
yAbsyi+3EP9JlKtLTasJv8LcmKGFoag/xlaalpfs6h93jyqBETZl8zK9vIoeX6RWUoNz3jlkRC+z
k+dAqyZzRkcr0lzh7juhL37pKoLbr0RSJzh3f+Bh22TENwdeFinsLaZR9IRn8i8EwLwWfccROZJZ
z9XgKz6ZhdQnFyZHL08542F5nC7NqZ1UJ/rpJLj9cwBm//G7O87dsd/ENieOVLW7XRaNX8fl4AsP
0i5a1flqy95+uW0J/QIpoHHS1xHNAZ3odhUs28RHmDfvUdzbyvYN/H7xZAGQKZQc8cfmft3m9Cx6
A2CsaQBVfNaCnxW88pVvnCEwVSR1EYZ+b2LQxVh2HQFrhFegyXuma3qCQNK/NyOuw02TlSPLYkkG
o6cw+d8wj5n2NJu+QX3b0D40n6RYhAduNrRbh9kGOYNqezK8BP/cIxVv3UeWWMWY2PClCv4gL5yc
NAWTJMSAednuSAYHat38mwYyR/seqFoSR9BPf22TE2LCGn7pJnUdbCjc26WryfZhIZX4zR1Kx92Z
bi8xCQhsqc/vqCQ3gL6r7g9p79NjR6m87rE60m9b6LEdHAA3iE7BSOOt0hUMsQWeTPC3ofh/e3mw
EzirX1YwGR3gxtUgM77znc0IKF1XXuSlLJbP9McyvwBkd5mh31Ce7pkhdOG3fRxz0JhVItoR7nqo
fQ6Yc1XdMaCKol0IzQqef4/mhFmDV/Mk0m0JZ0hespLQDLoDg1k6Ntlex1HMI+PVuc27Xiv4EU8t
GD8OpbBQ3oqjYzVcUTMezxu0zrIPmDG7BrRtI/4ybn2lCEfaA3NdS+QSMEAT3mwN7eoSYK4aSaPD
Nc3I31TinTE9Jl+ZGjhsqKT6SM19l9TpZGb+gVQs7Sg0w5A/6zMIOUXJ+L1WnF5WQQBttn/VX+QE
QCioeEu+Kf2BikQEIWBLLPqJQp7P5yaETl7VDHK8n0q5osmWoyD4N7PJbWkEoD7D1spJCRmiPUx6
1ol/xce3I3rYZHW4RaIipukd+GHrnq15rtYv3IFZ2zzA9EpWTtzoE3D91a9sb47xEK3Of43ZpwWw
fUOjk4DUjd6FqIB6mopTcM3OdYb1PD3tgJcM9gFWdtUVw6Vi63VbOhbxQcJzd07elM3iLqF2blWk
5ALyNGtIAiQwb1217fp2hCk7VwFMMbK7A1torG0FY/MTQkYLwDY6fiVkh/t0yUdC5z11f3odvUFr
D1QyYiyWobHexzqmyNEGJncZipndzcQ60u2Jx8P5/rvrRe8ytm+U/TfNiK365WubribzeVG+RPo7
+94umA5iuOkxzeLTjq6Vc6brp2R6l/ei4lDUtve5Ald08p30cTKhb0RZkohzdYIhBafbgnh1ndAP
dXC4f8ge+WLJKAeb9EMxQIcUr4bZPOweIrZTPDiX2s6MdSErpA+Lcuwfn0Qom0prJi9skQRlsJg9
m1/qk7euyMY29gvSgkFuCxjC7otkby5714j2mDYUE6yg6Z/HPmsyb0Og20w6tx7IswXhgfny33Ik
iCvPFETgWX3iAKVfiCARBtoBV2DybuJOX83xIjUObEzSxc+ZkrbW6DYiQNHuSXXy84xB5ertv/uF
zRvNRld1VuLVtGTrbbGOImuQOJRXMj12fC1IR5nN7/lhB09gy1fWsXZKwH5MhDg2xbZi7YNIKmId
1ZqzBhJGy+jdImBdrKAN9BrCoDuG1ja44BCGF13n6lt6gvRAOHDgxjmWv2Ag/hpjzagdDKCwPvP9
gzVcDClkKpvGcLhk0wVLf6GwHyjgTodFcx/zy6XL5M3iYVtGJyAClFkryPmU2JttBYA+vr8ZCYr6
X1icDN93apt7ldf3jsIq7iAWuUgj2v9w+sbMAwOk6yLXLTS0EBEXbQqPRhDig7Hkxe02zmYwk7d4
JMbtUgczNgXjhoBBIsGGdC9Arcl5oSc4DJ8MoBC09g5ox3CoWn+AqwAdcwREKR50VEJbjcSwC7UN
2TEV9ZrzifayyIvL7xLn2aYq9Q2PTR3AAK2gs9h/i2ywDq9guWD8Xp9FypdQdYwlvhykv/HcQkid
w3+L4JMAB0A9Fvi3EfAmzeDtFxEXgLNe6E96IaA8DwwaecE4Csoq71VankXWjZcubijFVsYflTcb
M/WrSIqI2rYkXSr3ACgdzkQKbhz9Lz3dG4t2FwdrdBHQuQ3BVgpbSahcnQHRnqLk3mAUd72SvGdD
rneX1jJCu/IJ/3zZNdAcU0LFNeAVHcQmijdRPIBo+313skDCe513RK0TYQF6Mvo6tArrzksR9ZfK
YPP6zceKj5X6QpQSI4z4qZwNRpJoIrV+ysgWO6KXZxCEqA48UqkDwUny2ncsA5MbQsd/1tzyplLS
1WK1fh2bXe+HvMQeyUXQ9ih44HBqENw5dzLpVXh3Qn4oSXiemr9NcdhKfDQlLD30MjQ7uAKWjvMf
F2VhOTh9++9PR2w0OLOLDVIrAlcodYoxALs6y1n2iZjZX0KYZSIXaSHgCeqS3DQ5MrQhFGo6L84C
77dAlo4JWJ4FXKw9HN5gzG96k22fN12uzlOG0vUH2NLB2v/5GAHnUDJWZMzxFEXgna20naRnvXbu
ltxkgvynFn9nnIBFQILNzQBH/8V5kR80187so37Y+8b0eAcTq+BM0cXiwi3G+7t4TJg7mAG8pTTu
vG+HsXz2j+IoWi7ZSUQlygv1UXwcylOghG1iZOh5ke4fjm3Yo9i6hDxGBGDJBiKvU+QgBmfRW12i
ZTmLqeFfyIUC9Y68Fk7/T5r6aAjIo/M5pfMnf2fso48UmCdWshFdbVsOz+l1G5fEXwv3LOqlW/bf
5lGrDX7fEaapdtwft3M52drhBDW18QmY57sBwEgmZd4nECL/tU/n9nB0nb3zWfOkWvEvUMeziqsd
2CkCRTmCo+sJ4VrWLVhgeyQIt1+LeJ+9/GQrwo5SWiZTor4sidnRUyyAGYSgtvndy0MeLClZ0Sle
VKJjKcd8NEI/wEAPLNbmEuELrnvSLapGhvTyjPaGnizeXbqNoI0RIKccjd8cJICOLa+ehkbb/p8V
QsMXxWbSGtuGA+s5nAaP2TfEIwiAjSNT5FFslAIz27pqiDbh4nvYjs5M0G8G9VsiaFgqjkU0Eiqo
p6Y8lQ4nLmIP4Wqds5Dsynax8A3JUwvikpdT5A4cNwxk+mBX06FZOhryFtfryjCWa7dvXXbkNOov
VpfslnUqYLWCajSBr0ua+/5jKuuyqZTTnPD5SrSwlSy9WSp+mBTRYzL+W5zWGWb1znXGosHXa2KV
aMVzIreMtUhZpu2rWKXwdb5of/j14hdv8HipvzA7g0Xr7KnngKhwGRWd1kRuYUoeou0UBjpbeb33
OoCwdx2D18H3Ipp4ECZp5IU0RnV2uH6h20mRYwTCLuM0BX/RSp6RVwijJGnkZvhhd4SlA/yJ2yPO
QCl5sxUrsTV1+4m2HST4dQJNGfwQuT902w8yWUz7QMdwslyRV0BZx19VLBNf7eqAQI/C7JTC7LUf
pRk23XSvlPIW6tlCD3e/7ugCEAdB2RmKPrQ0mhgZgHVa15TyhKq1PzHaKV3qn2B+g2ZU1sbjXV9z
+VY151oKffoLV7nvMZ9iVCn/njoNOFwSDHd74eFROFbTBjbGHNcqIn4HzXzpZ+HaKxjcKVT6VSX9
9Nb62j6toaFZavWwrdGN3lDeRUUfa1J7swycoTfnWySxxOS8BSMhXeO2u0SaSAN6LiPgjNbztoRw
7ZWgI6esdkUrRFdREhFm/axkmWU0OX8PnzSZDHaPsdxXA30HE8DacL7XkUwohRgaHNwMGYtHKInY
K9JnX3bFAy6UZAj0AmobLP9+Z2KlKS1DeW8K/lVLFTh5exPDi20vyBoYaF8pfJVCfVfClaEJiuu7
XKTM4tKDUbPfxRd59kQnOm7KeQHW3BKpfYuxAlzIyzp7GFsRc9RQnrEQGfLIFsbWGU+qtpJiMNR2
FMOE8VL73dnYPbYKUC6HnrNMHsL68tdITb2GYrzwMPfwOVhmHq4fCn0xfrvEEQ1P3ps6YsH+jpnS
OL1sraf9s0Dj3XcxO8fEfHFb0encqe86aIwAYhFSS6PAwoLZIPRG3XzuoHHv/2RHu2ZrAROf96L5
nz+/+MzJxcGfuvvU4SmjZ3bwpk2vqRe+oYmFNqs1GZopmFKWhxFnUEy6rWHpBRlhwi2+8hzvM3X8
jb7t9S5sIe5JRX2csHIc6d2EBSdqG/KCRbQ7IgPj5DuMrfLyy5Wnhs5cQbshbgdIf2b1VBqWurjF
JnMLzCFvLY/3Wz1KqV8hhKuhqcI7Bh9NwDGbaklePJzDgYux1XzgvUhCWnNk6DZSsHGUw8HE3HaF
f4s7U7WTLh0hQuGzjlnWm93Be3gRlWahCHR2H5BVi94pmatA9MCm7A5fzJIAUmsvMNFMjNOtsjWs
/ApyfosT7U8fl4NBwdLqc7gfAtjaBG+VUg+28jJdsREvHriryLdGEl4YX7J+GD9HW2kmmk28CdiI
dsC363vkVpv+T+2CZeTfSb6rrzboZQjyic7aqp8nhtfeIYw52NC857aCnETT9lSdl5PrRDj3mVrg
EK46zJnrGX/WfdDIdE65Ia9AgQZm1WoKzK4KxN5Kz4N0e4h5fgaha7+Mc8fJIHO4MYHbVWlIMLvM
Gtd1h/7tni2RB8FV4ak3oNSh/Z2opRSncOZ9g5MCk45jsKNpu5Eg3WkWls741Jafav7676ulRobI
V8ek+zDgBtZ5sxPBytHWIPBChQG8/mldwJF4sZGZE9lQyZq7ZiCrm6cuxiZxFGil1NjpA+Yyu8/w
n8IMIZESKweTdVHPgdXrqh5HCfU3etT2B50S4xe9Ao0d3B2kpJukSIHBeqcaTSNK3foX9TFHrH4k
03IFE4n50eUzWLBHqXkXWWxof8mdf+ONc6tTFqDyYH76W5+xUPy1eZ4zJpTQfqL+zghPGrHkUmtw
ra5cipcaoTNM768nOT2X9HB/saXeEN9D0dLkQA5HNnF1w/NNf6uagwuIpkt4ZD3amLBhP5fpOSve
iPU605weT7i+6G+TXhnPJhoikvBO9Q0cDsCjAqCMtA14jud2ncbJ8CE4PhOwiEyF2Xtp5QhylSDQ
1Ly9HAGf0i5r9RG60lIpQUCNgsqQk285/ST6SOAV4aJxk577b736fvqAFcKUWZl075J28z0wq4oP
/bj1nVuUvhlt5fgGM80GXFNPWKj9KjlP4liggpyQGM5E+ODSe8eQraXnapzN9Af2jaVLN99MPQ1T
BVZJOr6fisFQZmHu42PsykPluKNNIUF8w2VEssS9WoOftyAcJ8u8WB1E+Xd1/palqLsy24SHQ4wT
exaq0i/taXTmyC216Z9jp5HcsCApxxfiFQc4l7vLr3QYHp77u9rJ65zoygmDnYDgxGmK6eqmXkS9
y3hryWrjK/1C48qGrmUlaDTA5qZ/KzG129lmoh7x31Gdk+zVdG5lqNJmGDIfZFO57qbTl9TM5rUf
nFtbNb9w3vg7WUrXQ1fAaovVtfVxxa8q49n8ffw3qeRBOa+k/NfusrRUu1rUJISTHE4/zGdDR0f5
v/2lJGT8/bEM0UwlZx30qvITrKxxfAq85qNY/NlAQyI3tNKWx82yP+Jn3QVW50OUHIA/TNoEEz5n
v6dczBmMD5kvdbYPwH0fox1Rnyfj/UkInweaRVYGgli/LvP0I8z28sQDD1jWJw6AHMFjPg9Fm1aJ
tSlEAmVHFKpDwYMNVb9q83pxiM9XyZ3DcjVClYKnTiU5uICw59F0/mKo9frK63GPQlpwsINvBDRj
eiLnEGaY0Ltd28yxLN26OoVZC4+67UrB8W7aMopGH9+/Xor+zMgyAo0AR8YAN+6URXJs77i7PD2D
avOA8gHdh/iN/YZGL3N/OEUdLGXS/lGb/v3i28z5Hsg9CDUdCjWVJ6867cC6SKGSK6462KcmFA8d
WF42WP6vBvCZtkJSPpegmXJPWbRD+mT9CyJyAinbxfxW88rU88j7G4Vi050e1ySRWO6iCvpsuV2i
VoS7WVSxWti0VDJW1PVNivibCoO7Vv6E/E4rKdQ9JjnRHiCjyjeXLLglfZ1HQmqrHu213fZYN6PX
YFWyoait0t+DWAvNF/7ftCFxgN3otJJYUignq+uUQt8uIexT364s3bswNeURIWnoL0NrGgCN+hpb
6Nznaa9jjwGBNVl3xYTi/Ic3HoVHVCJxVswcq6X6gKmPgmWgLBQkTn2a/xq+qRLPQ1sqL658thEa
fLJ3JjS/71LlJfzI8iokxaXl6YRT6dBQEy0uwxanSkMNIOLyZZ4upcvkcgtfXhNlXcbUavAui8f5
FyM1HDCgNIoSZ5FyjG2LWvzz+80uG2nPeNJR8fPE7/0zqE7Oq2bdWViey9LuRNW3QB5p3ySasOUA
OaJPu/RQbVrlJVzyE1HRuMMiebMnzPJ5NZ36sukTLcs5HGc11uyECTVVIbt0Zu/z0gs9/zDzlhwF
TRcm14BVyc5aJAsTUUobNMM32+2Q/EDj2lYLhdNFEOqEA8scMUWl/Xwfi06qsmovSaZRsps1MjZ6
rfW3iekrmwIdxdUhIUti8rSJXrzXzRHvf7cPkI7Zkx8faqJ3YZTXvANP0v4N1xle/gZ2e7UuaGUz
+5aqvj3v4I11n6I9CU5VghQ+T313kq8Teh60OD04lJ/xCrZm9rUVKIAXpJoVSFA0alvpq8pNyBzY
dTd3PinRlTM83hSiuzgeT/qrcSJW4MdtlRiK8ZO1GyZ1eZVU1fZZttjvL6DxHYIQy0pTo2Mqc2Oq
j5sGx4fdGpuL/fsH0oRLgrLzGioIc5nXyD09Z66aMjOHuKpsmH/tB7OF7/YCSfm/qR4tgzkvpwLT
5VWBSe/lOoQGwK9Lf0ybZDpMejTWUUQC+XONPddx4GkyP+ZKOvxU9kfyaoXAcFFukRR3qQWU33U0
PaaHLxOEEJBTR/3/78jv4nVV23kdt8qTfvI3AvnLFULTNfxsl4c4QaZ5r/oMDGxB8ETGxFDK5SYC
X+RxN1RVxXxxjiuZzRW7xbXlKIm14GQ3qvuT4A+AB5adrZbyqe9+V/sQYgZnYRuzsgmIR199Sf76
KttKotQFOPQC5nSTsjtC3ryCvPhmDxiV7lrJeWMA7ulI7I4lly8rwxITjIkzpo3SSajbGnv5MJP0
e8p8th0Yg6CSPOKD2lyIMeSDx19tyL2ruRaTsfNPcpqWu345KwFYpRVWRUUL94akeKWhpycSI39O
N1zMJanrQpJ3yBsdFWlpTNZq3KwsWvNZJngPX/wFl1dAXpwiCMLPD43vo5QSFqrrUlj0Z0u9BFar
NxLo4fMdTOU6R0HowK8L9ereVQUBdJcB1UWQ9RqR+QahYYCWiKLNVZcdoC+MWjZS+opuRtMFIINq
7ue6E01TZl6cdg3BhK6biQ24iph6fqshuc+NqMxHGg/6YVjb2qXWuEMOVq7e4RqYKhzSxOKQsOuJ
3uv6ihLVc3XoYnemmjgP8fVbET3PCno97/FuiuhwSyA8RPjdtINAUbjL2a2TX2M9sCBN4sQWJDLZ
ahYaiSq/cJDrmj1gR+czJ0mCE0ztE9cgRkpJLmqiAYx50usnFLapF45WA6J4WfmfUddSqIjfg3kg
BPgf7oAPOLv34Nz0jMJVv9Klc8QQ3+WardrvnwbhT0UXASPyCOvyc4TOo0tEITlp9H+9Q0HaHoup
rPA+QZBbdb9Ew7Q95d6w3q4U6JXESBRI2ANim5HrXtSIDeamJvpojYvjFOyUU/kAzXNSRKli4zRJ
Qj3FErjQ2yfEFYgU7f0jF5ii3FCDpacFRxr8c3Gi0sL19PnfMPrrVjm3jZHBeKrIHnVZPi2rnQ/i
FmqgRvjFQM9OKm//RZzQrttsvDwW5S1bE6GFzrpu7Kc2eRJYH6t/pS9PHMIle72jOsTZ3+wJz11C
q5+NhdHb/xxGbzYm5CZXYbEjJZPiW+7ukNe3SwyT4E0PvW+eNDJqEkbaku5EUIAOtwthmqqVWO9V
5ll/SBEZq1UwtlaIaabBx76mbQun3NFC2rrrGaJodJaEFax9QPZnvF0hvPaRPz1cWs+BnrrcD8GP
CSzOkPjfmC0KxN1GqEkOb6dOCxNVE43uCZKS7O4Y/6GgC/sI+qDdLoeEPDs/YKKUOLPuBAmxbgDL
cCYUWme/NZ72Z4Ngj1MuBXsqscQPY24Dj2KdAUIBMrFo9z+OXdJk0chgz+PlbvER51SoFk7xbPwe
jUeYYspSI5AueV4pDEJZ6JZSnJNaEJP4QBm2nf8isME/ooJnyBFwtQU3/X+WvBsfgA+3BGliP3gx
7TDSdFGDtAtVZFanGyf1W0lqdZq+mz98h1PxWFr5KW15bsAt0U0Y5QCUO85CZnMBZOc/Lrdy7+uI
kxsF3oV/1HuaCWa+cVNyhKCwmxMKUHuG6vLTVTKiwhVlZsu2krLJ024xpBq88YoHTlW7Ah3nxe6j
LmF+bCMiMYpPDoCT7+sDOlw0mIv9RoYw1CfFfynXJIoh/6oC02ZD+jv4DKqy4eccsIN92IlUPk6n
YIgZ+km8jxBLfj0vVW/yY4PCKdSV0mGR98QvtAFJD3mCL0/lA5ExCLt87fGwopQ2N1fJJ9BWjlxu
nDxTX+EIHJkDAve8/Up6uDIVt311TccF8+Ix74KfPN74xqE7hRdwLEYWkxN7+xTApQme4m6W8xxW
NVyHCDu5cwDXU9V55xs4YAjl8FCcPpPFVbP/mcNOB7m/sH11vAeyWgNl1zkr4nPL3oCpw4p5f6XH
pTbjvOHYdEeGXvjK8sV/+zVL5yKPZVVSG23tmJH+lfKAGX+BTGhX6IMRSMHtlXTpo/4XfHGwP2bV
yrZlPajI29DF3/oaG8YueJTacbRMh93J5At4RcAmloQ7lk9jYU/kCfLgHCroREH2cO2dzt4hcYQ5
3H9ByU30Vt9NQVll80X2nEYYoYCAOgvLRTtj1YahMQi4h2Hf5YUn68t1InXdbiuveF8LWbO6gDPu
lP8kNEFT0N2SFIL/lLOcfihiFuBdKBsL5mONmGQQ8XI/oO/SDI8iNiftDLrlDsvxgJY3QyjaRCJL
JTfsoHeGXp+LsgevF4mPQdw6h5log9MEkV5Ky01crMFXvmX/LuPBx1F6EcGybepMsY68SrMXwVMR
YIavODv+9ELIZXPod955R7lzvzB6wwhb2U6joCWhBDPwR562Oi3YyN0NK7nxh8EpHiR/vPgOa/PW
sg8Qx78+AKua0aJzf3UoZ6qTYZRV8LoD0aEg+2mf2D2fhuHAzTtkp/eAJVuD2KXsHiPrLGXy0vVG
IeCBr9ztUmMLZQ1+KWojEkH7ubfBjLQ4j4BNRIoTwglucbBKmzuVb29X5yuQ4HAF7dv5H21WBpzu
Z2dOmJOxNEzoBWmhi/WHOmiVcrtKrx+JUvv31zMkz5UE/0SovnSnNfm7a9klBz2Pq8fVP2xRVm8T
NdfT2TlJ9g3hoF3OvbK7SYNMxdvHW7yce3b4bTWywiDvnOPAP/mjyXg9xFzW0s3RqMG4hfT9ciiU
cDce0qpI82+Ay+J8mHmPf4RiGGQ62dejvZilDY2XFW1zjoUS8If5Tx/Y/6lB3BUkUNI17jRRuAK2
q3Q+wHbgbHWwFvinZ/ZMxffLwd6X7tCZIFWgQTWcJMNu/Cq1s78rm1jO/W/NwyzXYpfbJPCSmzYW
wSt5xqFFPGIaQn4ySWxbeyngZyT3sClpl9gnM3RQPUfU6uMS4+ZA6US6MSPWtkuuFAe9oN3G784t
PviinMKUohqCWFpRdCiN5miAsu5Op20oqG/GJtCXk3nn21zU6cS7ZtMH8wdaJintj0/hLsQuNfvZ
0aMkH5hZgCXfWtzI7EKUCirkOcEQ5J2KvB7KZAUPWJVtA5Wk/WRcZNAqyd9eLLrD6QJ7Ka+FXb7t
hucS3FL9ZjLmZQ7ATiiJ5AQLrcXxhp+Odkbvm8r/lPLe/P7EHrl4gp3MNB4lKxpCAVYcnGVKuIE6
s4Tuokzsk5NpNigzd4NUZkePCdHK/4668ST74n1ghl8q9L/toOih0gIuKY/vebXVqVxQWyXsTS2C
w9g9FR+pv2Sfj4D2XsCbzqOJrbVhazQ6KaYnFb8olosvrO+QGv/lwxh9HT0zqsYAbLHVwQxHjeSC
UhvwVRuJ3frPeDbNnrx1QiJO04n91iY2J1KHe9DzA12AJrzbo1SeN/u3xnGgg9KWAxD1ZN/FgG3r
Foj5mr4HKLjrYB/YPRYEL+vDsXkivLasTzMtswhAMrRLCEWs9Hfo14iyaTm0+a4ZQigfKy2XvJrO
o1ndt41Gcgqm++5w2pdjpiwsYYgRNfzFxFeaJFoS34thGiC6u+P0EW7/m4TRxdDsu5mBetppcfqL
UUNoGVXevyAyX4hhIdqLXwX90mn5ZokR3Kt1yp7/edzxhxfocx8rq7P5WvaQp521jv0YmBJKXvF0
qrLNqFurSbA5N6mHTr1AYoaT2u96Uuay3W1Wk+fPwu+FkYpPX3mu7IrwOX+3BeUYsA1JCCvzAS4O
V5GILRuZ65y2b+GvyME2Fibg7iaEuDaaWMF6HJkgDtAXfHjxVUq7g0CZvgiZDwsO3lQk7ItXsWqG
dhnPDHaqoqe/kt1myc18D9kJ6Ag7+uIlmCe/jq9G57wk2bPSECqdytyKhr7vXgyIlKHNK104yNAW
QKIdMmw19C7PG9ZqrkioeXcWBCdK39T2L3lUszWYVvKdM9TbtFapPvuq+axyZblS0fVnGvC5b60S
/4oML2chRjBItjEqT70gb/3C2Kyq0L5zlrmLpCSkhqlBa0+1yNJ+fi3n37CBMCHvxHPpvZMvq+s3
RAqT1l0c2UxO0U4lkFUKUL7uL41xwKBhuY+RDUWilsJw/hm1Z/ixfaLdydCHSYJ26oYPD7LPRQih
yrgQMek1LSF+PjxT3osYIWtJsesJluvF3Vevd2h+p9HWVQH+jN1mMQ4HN7+5SyDXOxL8pvf/Icrt
l9TJjTGgQIIQHb5Y2gKZaIUcZSxmfr4AWhvneV8VRWQ9+IDRXITQcqhuME7nwMMYXt3WNgatTcLf
XxbRZrlEu5X67wUUsos7JlWtpvMqhU+nTJsFihx/4a02Bik4Y33ZQbkEjWahKKLd1yOnzqAheaTH
0LDEPnisso3pnD2cR5nLVxQ6Mc3Q1mOqBwHsYZ6YDCjderYIYDAYc5UBa3wsFNKUiW512clXec4y
KoQYAnHhY7wcc+ztw9+1u3RU2YqkMGJ9tWHRVPwY4NFgA3GkFbn4j4OTwUURLu+C2rLEGgB98j9Z
MFbHLtvGm7Nj45zIuXNofUFqV4AqYIzN82oj5yBXrx2YW3PmdaX90x8n43l3CsNlZ07gyCACvMA/
rxb9niJBfOw8St0tZYiK6BukX/dKN2XmXvsDYwjIOaStw/re9SzkZpJdQyLlX40BJO1Q+KsPqKG4
2kW3eIVdl05JlNmExaCyeA9mzLl+T/qw8RPN+V24lxWclxeh1WRAT2uB8RfGhJJydfY70vDImiJU
8rlb7hNFGjFvwqnWUz9Zd5+seLJpE1Az32zR7P/q+75rbZ+W/wC7ljKIDvIMDYNeGLLRfJZGKcxA
E4eJQP4j79lhmUk+BKvjsy8+jIyQMkV7ZWT6Yy4jD54BJY2vfuJJQO1QBefbaDj59IR3qGeF4s9X
6OtwzEytwVev3fk2l3O0p039Opm/mxaYjV00Ls6MOuOWw2RLJOFULxcMPUgyiytyXmmJOTK/+fbC
qkYQUydw3Ip1+JS/F90baGtmLEDZwxa07H3J9kveAnFFj6Vukt6TQB2VADS+HdQ0QLFX6TaUAekh
ZkwD/GcmDS++CL8Rvxry7KcGRLLufceqDPUXFjgJatbM3F+iFycOOc6SqEubo2yKCf+g4M/PoKnB
rD1MZzmt1pZt2J2zYotbHMo9URd8i5XUypnkSJpkrPWRJcyVsf64RkmKkEnLirVdpuTc/4kM4U13
M6vXI9Ezt888JXLAEUXPpNN44+ygknYJMY0KREUnk07nkcNciM0FtJcdSt/4eALWWcgxB2MDT1hv
c54WFaf9LbAQ3T8Cx2kFRYMOMQYPfoNOTi7JNvWvz4wM08Nb/i8ee5V5LnDPpXvIuhU4g6so33+z
7LAyL+Sl9pp+M/RRIQP6aAZ8+dyTmrhFPIz3GKSPeNbmtcQdvwwv/ltpXGWuYj7dKDySTE2F5cfI
Ns9E5uxLfLoaId1OmKaA1Sym3zMNid2V37LjDdTyGBusiE2y1YlY96iFOisUvECKmjQVd39wlMBs
IRAPwqp0haCTGh2/Qdy98KDiUAzm6V6ckDiCMgSEOKsCjYR1oLjzqEjHQHuGxRVysFISA17rKNi0
0exC9JBBXVVuRGHzXTnWDwZIpTp386YuPwcSFI7wiuR8DOLaVSaLFECwMET90PH6RF321DjOCD45
p52IlSURK0BodeXfq2qosgQJl/qBi6QLLGeT+2fRdxwwe8okAQYWuQ4bKuJpYabGqrGRrVtoYbSj
0fSoXA2UrQur4XE2fcwfVGGiaz7TE1xBXOzLNDaKN9ctYWtkmW+1L5ar+CX/Iwt33RuXNJF1XIzL
8MNFrGSG2U60WaRiePUWpNndhOT53EASjTRQ57ahfFrUr9kbetoXXmlUyhiJv/upy8P7r869zuHD
GYqzJNZz5XGoosNgg8UbyG6T6j3fEpGN1Tuf9Zbit/eQRGp6dMItk4aiSzQ6iLF8mq/DwzLJqQyy
X3Gh8FOLABDGpu37Ellj0+qb17U4P2QUZundtwJrisiAu6E2/p9OT5/ghRdb3epcH5Nqg5yms7+y
OYuL1bjh4jYefig2NLWGuA==
`protect end_protected
