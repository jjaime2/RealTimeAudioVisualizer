-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oHHrCbtuzICtrHYICJy8X5NynPnE8v2dS9Sh3cp0WD5kyz20LmCmFj0H40sBmBidIybtsDIjYhEb
abTG50UUwQTQSjJQJ/7NBEHwXXOBExs2BWTtwF90G70YEEpSDEdyaXjJiqLZCqnqzrmatp1gutbE
li7aXo32tlYpu3dH53eN8sq9+QV4BQj+OolvWXbNCbZJMZZRICTSnkhV6d3eeQHXaf9flEpOR04T
qWLSwHXpnoiHycfKfMo+NLV1KCJ5ILoeG8FXsY4tHv+V5yXtyDQH/8ypM6JAUsfB2w/yUNbEQ7Ra
Fnfrs3T9Vfs59KHW45r8npcteBw9PuVLr8UJXw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6160)
`protect data_block
Y1z9Bb5S1UjpidThgtJPYgNuG+llnVHdVshBjgD4zy+5ikv7Kx5K6Y/xwWqLtUuCJM5GzMusBBWy
hsoDCXOMhROEnIhTgOQCHGqncaUuSibQP1FXbuWKh8yquoLgbse6Eq4ZGYtcHCgiTMqfubv74qqi
gdRQUBrapfoNbh1sCvPykB7c0JsG9J2qKz+nY+VA05t0ceB7N30DSmZ03UqHbLmjBZEnHk69S2yg
cmUDOfpYO9g0j6SZpRC+ytleaEPqCoHOYfGvgP62/2lXBcJq6/l5H39gZ2pn74NnHtCN2JEZpkwi
djzkHwO0uVZUzDiig+rKKrYnzSNDJwvcIc9YrNg6yLhr0vCyTIDX/FUuQfZhjynQHxpXou24uDYM
fsICkRvve4NnjxWJ5KJNup/olXKduJxjIn5J8Dt5iVNE5jS6IsYOOCWLiMkhyYNi2MfnW0/lZfms
bLVd8N2wrvGLyKgvqMrai7tSdRU6Y8lopLmVg4H+hdTZPRg0JFUvMrzJpE4j63Wf9g+zCdZbcxS7
fjklGY1uYc/oTZGRdv/jOeUE0xPfUX76QjK4bifX2keeDOxljAd6k3Na6OVXSJMEqA3W8UkMJeAA
tZ6F4ox4FZqRScRk0UN5/34Hth11fIIy4EvXEB6naBt2BXEMibrY2lsfL5h0fmkUl+oO4nMBIyFd
nCBwmnGfbFYFu8YJaoVryc6TeUCwHSmfD+tBHLXbmeXLyu9ZAQ0o64uK5vwITk4MQtUHFOLq7Wae
Wbzk6RU4XqWh4L6/04JexuTbjUxGUbjWmQ8sHRvgeHCX772+Mu42A6acDTUR+TiDkF5HX7sj4WJ0
R6C2TMaUHGSMP3uhs3hO3ywUPQ6QlEyCMzCr+xfG9Y0Go0JsQDBzTA948qP5KlFJ2dRo1pRIgvAX
VaTMxVn1SO683mGHpeVce0dTJslSDxPvbx0egBA49g0fHRkcRY7pqYuTAWYYpp4aZqRWL1ERMm1K
xywx/H5CsEjKlAeRbeEkGLaclyGu/8MfPQQ80lth4EklGoyyHPC53r0d48oV9qFSkk8Z9zv20OXU
QVyxKtpKx1BNwYirbVCKV3xw3K7tlb/TgtZNH5UOGiolSnFByqyYndQhSMRf71fgknlUrAe8p11M
3mhc+fx/qfSuZ5tNVo0/9+K4o8fPOntchSiJ+i6iSm9a2u/1/fkZprcCxpp1aeSEllspbIH3t6+c
Hg/EVAtF2GXb/0fHLEcLOdZKmNQi62O2IsL6yvhLfJcYyZ8WKCG2TJ2XoM0kJL0p93FwI1Di1CJ4
s5TQ3155+t2OIvMDBJnt1xn7SXRS86wLYEsbIfFhQ6YAHrQXQ/gGlcn7mf5FokM8+7eVhPYOQ8zr
DGdSGu0+/NSJB9E1BBmV6W/i5qTc1vLWxdAFiesai98ZSEM+kW3D2cWP3Pn4jX9DLsvVqdWO4q/r
xkg8cvaB+bebimPsE2RMXmgRhByu74uXQ7KgqUqIe4gw6xTY1Ov0KM2H6Zdn07ptum1BoJqw2OP3
5IRv8Pt41bvW83v75aV4nbxvxhyfLtkBrt140ZDyIQk1s/Ti5mtL01RBABF8cRGTRv/uh0fPpFvH
ywHqBYikTdqXJMd3BJLY2hAJ2ri1+AsNE6mOuL4CfdwsCHqB6hI465KB+Yxb/PzDAboyipNCuIsS
vngomfqPSTnbvwoco7TmCY0y1+PIc4H3eErnQtmV891utav3sknWgx4OFpQ5PzB+aPSgMZZV1nqA
FN1Vp0zoufNh7Wsp/3vQUolK4AXeI7fyV2pgLJTvyN/F8J1XyuaSGeKIoB2qvMGNU9fWBcM4ehaT
XIX7vuQO8LuoL0ttMWgiISTKpioLS5R9j/5SiRM0d0yUqsOq2w5odD6E4b/RSp6lmnexbg6jd9Hz
rP2Hr5kHt2pbiZu1OPJ5PRxfBiPYH6naIMXrTOxDPxw4gl06wqK83xhSVtqVhHiIe2z6HP6DSFJI
NTqfKPB3ciMgxlnXzfuFVaFV7A4lPTiWOUFcgYpD+NO0Yz40nkf6cluMOHZGs11Zs0uEiQ3JINXJ
fZLJnUelI/8QF2I89JDXc8mE0cZM2eipOtT60CzX4N/c5zNUdSnYy7Y1UOMbQEmqdjlTrRr2kVnM
YtMn+43JI6aIPzecjmMEWMjXG95dJ7Ht0tFNYZtEm1DgU84UFwD90N+FUqR+he45YyAEDYEIQQZj
Biz3sCd53AyR+TrWZ8PyGYHnrEDV/gyAG9sTdadoU9okF+Vboxzc2OJ8INXK1Il9BM2nl73Mw2Gb
zkN3W+rm/2Zyt0Ivmn2Pn41+L7VppHJMefCTKgjWTAKs1kvRb8qhnx2QZFWlF9AF2AQ9iuXl6P6K
t1EgskmeMjIREiMENoDkm2S7p+HY/iSsdrmqpgnvsZ8Zgvmd592r/RV7rVipPRwZ3c4jqh+6lfRZ
RmHsgtUDlZUda5mFBBdd7V3TV8nlr+3zDvye9IdYd5UMb58cH7C4ET/7+3N/InqREzK3FmBggp/u
S5AG3tFMltBQ8aO3LLHN0st0oqxDDaEfll0kEjuSG0+Ctrw6QYpHLAoG/vMzPQCHdroRN9dCuNW0
+Z8PWSJiQHzURm2cG2YJIZTVGjIUSc6VqXk45zkA+cFub7hlhxAz1iV54nYFVFUxYnA/9qK3jIk7
A8g7dtT4ASTbRdzB8jky/RCGJnrYuSHKNGQZGQ61RiZmM2OsvlSJs0rFmln0nNAXbC5UEjAydIy4
gsPI2YXouDe4Qvm9zOmHKU0c9opMrGeaZ50hN8GZBcUnEACvysyFc3ZUe229AnlM823ihiM+dmtA
HZVEU31TcyEGMPQwLMeiF4ekRwsLrH07kcvXi9B4hanqTbjNRhwI2uP58leAQY+WJw+dsSdxnIEZ
K+yKxarVgIyL3eDw4I47vnlsy5i3uSBcxAZJWfmpQd7+/srO5lhxG1gQ8TcG9+6g+YrhPPQVtV2+
mx0Mzurf7lR3F8Gl+Axq2XINp/BmmhexjoB5hSYICfoc+c75yI4o24nBuDDvf8a58Mjfqc4+hUjD
j9Rv8Jbsl8sHcj7Opi7DW7WRYovPLzQBUsA6bQ8Or2LfLM4vWimi2v1GrTrvgBsHd5JHqkWE2puF
fUriUEwF3rBx8nS9ugmrBqncwRr2npoIPnE5cKe/j/84jowoBjkmCo7QIQkrSuacJWjCWIdM5q2V
l71XT/eyNx4feyvTSQXpSkenUcguaZpo8QsSNODS2nI/GEsfpDrDKhIMo9NhRapnlmGJtNftQqks
1oQP9nsWiux2ir2tJJyEZzN0YeisQCsBv8En6I9XuXAWKLiSI6q4rCBgX/k+NZt73eeBTFw8q/Dg
2aKEbPtxzPxHnDLmXz/TikH+8oK7WeNeADwTkSsWfWw/ggB2euejrhSik2D9g0rIAf+j+1JWd1xo
Eh4KdqL6vTWg8KKOaxLFmtqV+ssJpia769DUJTUxIlXnFEk5NUTllHeJ3olqYVb7T9hRePyPKkeM
QkWPYHKuQQGyjXzRQbUvfN2iQ9Ojb1miLlwFG1zU5lnzsjvisCuwBweaEmJEfSDkKl+ERDhKZe9V
TramMuWtXhW3Fqpfe+Q+OXKSSz1QT5m18rOorOumlRne+oCnmA2JoDtVb/Upw7QXNHhyF3JcJzFo
h4dPeU/wsGDgV37boHoNFJSxjMt1eKBLhZcUo4+7JjB7sLdWhK+zpR/LaA0nKfaDC5PMxQS4sGPO
d1yockanm1GOTs3jfZpDLEe6dhl20kkgcTWwKInN1OOiLzCYRXWv4tNE6tHAJOfXWSRtagCXF3mG
Llq5MS5EsKPnv8WTpg/cQoj9PAV12xnkQf10gggfYSoIUBgOk3Po/9171uTdaqWwYXH+j/Hc2Qq7
P7/YcfDeaGXnnmFTLwjsoDvngav4Yt63MyWb58IeYUNRm+cUL2YF1oKDjiwphQuELMiVQY3Hm/Eg
ywM4t8MISYmPI7OnFYZ/fbh2P5lN6izPIlI7OhWa6yNyHhnXSzIttd+FQyFwFaZHqpxP7UYhXdMR
TcmvTfW1irdxNObOCLlU42kcwPSXqtIdxourlz4T5H5kqx/v/EqnXF47rppJA9gUwFYqx7iNLTGF
bjOjAPWNS5tvvpqBmepJjSJlZzctHg7F6EJz4qO9cXLQkayfRqIbvhXFhBya/KeSkP41mIrHKfUr
zfzPocHyHmAxsH2c+zSptXvn2c7rhmK7xj6EKIHVaX064jDIbGIxtaKodHTBFzM/ikKaxB7fEwTK
g4C2dU8Q8MF3tS0etfOlOw8pc+p1OHhaJzL/53wbVHWNpGAHL3qwqg8Lwj0Geiuj3HAXjLAwllaP
9/2aqGqHzV/prL8D4NFkA+BZ7TXMqK1QX6npt69kMZMaupE2i6SuIj7QkM7/mVeKQ/CxMTddwE9f
Lr6aa43zs4KmL3rwWm654X6FZhQJLcolzk1pm3R3wN5WZA8DnLzKYHjKUnIr1S83CKzWCThBks/l
8b0rIsKax2ypScyPb+uy3RO0R2t0YVLWzAhKoot6G+9wnNo+nhJSqytnsDEqUdVMjjMO07dEA43j
hSMI/qqNhsvtmal6qrbb1We20aHXvDw5cRgQOiAXwuvog1Q0gAVLiFsIxr3V/kmwH57liTLmn46S
9yWE+kr4Aif++7GgN39bafaci94Tg4Hcxgo48Cdf6t8OpQZosIGkKg1PKvTXHwGZ+r2Y7It5v3z4
HA3fR/bqE+DUHhII+v2lWX4kZfccd37aRfrPHhFRg+7XKci5Ak6Q3+2fq1S4RHUB9zYZoxHKxtYa
Kllbals6zu16cAePN9Khwkg2eNVtoBae5Gq+04+/DHnUVGkgh4za3vTd/RLj9Y6JWninFYFy7gwG
uf5a1yNWtdUe2k0SagQ7gzU6KniJ49VRBnebK50CbHL66EZuxL1X5K6xiUBYDVg0RiyD6drnwUmE
mMdsvscosru1I2ORiGWQGhczgyJKJo9MX1ZHIq/6QTcapMEx/Qn7ZzoncowS+dG6AUTgaIc7It7l
V8TwT1ThlMsYqxnZ5dXKpqyaEum5+i1AXi9O38haDFnLDeUAwXZ5spDnFmVFwCa4Y61fpyoDNCTE
94JVHc0YhzdwA6oV1SPDaXRL3j+v4vrKnqvny9sa4hQhIg2COFiPaTj94DGaMmjcYsyavYMSFk1y
IClAiwjav1VY5yp+lAUL6ftgcFJ0lINcu+DwcPKw3xAuXgAJ6jvcw2OW82H711Yj/h0QXrbCFwje
2dsfdHzTQtaWlwqocPhY5pZHMFSDbddb4FVtHKFRuuYDTS1zwh/GbR3wZ9GVNQpfVZ5uUtZnJBgX
Z4V6xAWq0GzwFDcRhvx+0dxlK5Uo4FD6hlmnm0BBgiboeanI2C78d7MVyy0qoNBTKjWULVuAMIh1
VbOaCUYgHdiM/B8N4HRbmE1SmPbbA1Oai/gGyxcn8W4TWFuKXSXpHPomq5CtbK9bSC8YaERErrT0
0U7hOHJdqCM/PAHmTaWilgUgbbbHE7pbh6RFz7e3LhKDkatvqiwkFKsvjhqh+nPpuD3/3E/T0h2W
IsRDzLew2qrEp5bPfIsXkHgcGXwedXfQ1/G9oFcLuRn1G2HEiyCQYxbLfLSJLEvJL4pIm876LpqE
46umRTQe5NgJ9cvsbRcGdGQSTxin4JmYUYkrnnUjs9Ltly6vOfvQr/BssSjdd4KpujJewySDy6SS
xWxkD1fqlRGweG2rPeYB59KDwY3U7HTp5gyV1jYGjAUbAqc0lFc+uYjUaYRhZbG4IyyaBohNC8zZ
sUh4IPoKDmuVpCpX9mYVw+gqnyeLNuV6rfzWFO7biLwx64IFCjNW+1mw1Hz9XURA2icbUQ9raHIz
YecatN7lo2ZP+IUrn6/gnD07/QyO0s3Tq1fx9eGQicWTNcT1OLhpapk2L8IG5OJpnUqU+0Fmai5Q
UvmaCU/omejzFf/LOWUQIo8kWabAyblnaGXsMDLEHQUfKFtjpRGJiyzxPKRAd7VhtXWdUAlro9At
aYrJxWc9tYyA1Go2WkS1dono+dGQPqDa+vtgscCevMJf2jFnH5KuJKpFEJB7TbdFQDOurt4Pcxdp
a9kpb4k5oOlFsUIo8Kv6Dtdvw5ngi+umndRHdeht8hoBvBQz+D/tXwjebQ93M6f/XzO4jkBLtwD7
7+QjDE/7yMnFcznwFCYLgf1cmS6QERwlz9OBD9xVz0yNd1x/+aVAB7Q4RqJTTSzKllYuwTsQOiSw
XqUUiRF0fPJUuRQMpOQ0gUKsYGCOBzvjAP3gaVaqU1lrxmkmjuwk7mKB5iir9SxWf3ns6G4ysoIq
SMXSQSQYOhj3Vu/HrcZ2RDxLPwQamjnsNhFritpnGO37vi6d763CH4hk51VkdCP0PKp7/BunhHN5
zMCJ89tt2TJb59ErQBQZ2cTFM0w6l9U9VVrD61wmBlPyyS5TFJ+oUd6EIztWHUpj+vnTbGwE9Ay3
kByJaL4/594FmcaFf51/ORi17QO954TJ5fNsDMZqvD3xyQ9C70uMFHHh03b4nBqPmvprycwb54w5
BdqPSwTA2NykxzK1wCO4ZKUA+mAm/qlzPxIwYCONHxQBd9YU9HJTwXN/AUe9E3hADnQuN9aZU5HR
lER7bHMc2yTd0S4mdOIN/xNDj7G2n7SDd0+6Pgh/ZmMifxxbfEV8uGWgTy1u+Arck3OyjtKGHTQq
yqtmJfoW6+tZng/JUrsHqmBhzRB+4EgIWfEv2h35vahdnem6pmniZFCOYF6uEvtk+dZBTGnbpEEW
9TZLuHr6sPq+lXFaqvnq16U+7CRYgJQmSV5X+L03LYjTVm9z9WLGFdNb1AOoi6S24KmY1qdtLo2+
+9qpYuBcsaVDt++OXPX1hVbhxfnSyRY69p0gfqpljdDZ38TWMok3MbMGLx5EaXENGdV4wFdO9wHe
5486t76aJXZr/vOk1Oqyg0N0wMudO7x8HtvPp0dCh2SYpnW/vfwm3wQvsRtvQuatjckSWNGyA/Tq
EqZXgyLx1TBCOCLfK7MT0SC+L45Aippu5HB2ZkRmNULNslJMskQQHzRc2pHe1whn+pBO9XkuXYZ+
FUDU6Yyu3ifNhoZS1PMioniZRf5y/iBcRlYHcmMWTjSBHu+YBufLMdU8ecr9fu4morER2qCFsV34
OdKCt0hghqeiU9FJjDHNzFYx93Pb5YkkBYjMr56IIsdGbv3j2NXtWka3O5gCnaeUYbpbrU/TC78q
jdLY+CrCgt+0+79VHbvXcIHvTrUPfsg0EFzg4ScItMfEC1aSXYa4hEoXHFkvhNjZYYpC/uPwTF56
OUBFaNYpC66al0xscp+CjYTL91vE2CdFvqf7wHXMF7TIM6hOzCG6v05MmzUsPn9Lfj7beGXBP7jJ
l4AjcYjlEhQKI/IwklPXztPnTLZtQDDyp6+Q4Sz7qpnz7ExHXkFvEXd1ohb/c1XVk1fkgPZ9foRD
RkMOqkxtJyYHSH+aNRx1+UNcsCyiSKxjLU6IDl+MWB2Frbpc5UHAddStu9vzUPaPd8OmyMi+bogZ
XegiiP5Lbi6QjIkNBiGGc4h7iur5ICDLf9YXnh22PMbMz7Lk+fNgDUuQt5ELgqeMxpJ6rEwLmr+U
TMAjLSlm+TkAoLz7BUlxInNrJmEtU3kxzKlkd3BaQxtVzmV7eSsntRJ2dRaRJbPA1x0VhPzYmj4D
LTLRaTRsYGWOfk/7/oTJgvmhobRb5LYPxDYr9TjWZdKYleGQz1XLjBIg9DoK0NPiejbZlh9lSChq
TYKZmFaFN6O1gi6fSSxySy1JNp3YNYDr0ZgHNMonWdfS9l95m1lPobjEB1RMyVqg6OmPn9Jzz8Eq
+dgBSkrc2YVwvn/1PNn/Gbsu51UUVagzwlI/G+8ciSTGl8Fxw3ZZ/PTJtw1TlUTN33aD+elLvZBe
yWAC4X/A5EP6ht1KTpqfSsott7AYR2z8YCLttFCXMlhP1hEpZBTXNfoPP+cQG702B3OXeSOOdmm6
9RX2WDFS1a0XfHT2fPletkAbdiOa8KeN5cutLoYxYd5Acn/A7Ozj1MVugnJQoy3kjgVZ15gO1Ts+
dG1d6T+NZK0RbW4wIbYBTyLCP9sjINNztz2+ruxGiRXJKHGuHcVp4fFXpnw0MhHuXCSIBqm3gEiW
P9W8gjAPYv5ovcIx6aQcQGQMmVybk7P1uzfxCnAraD7rTIKReP9zHmcQFIKn9KwYrPUBVg2HsnNq
O7wXLg==
`protect end_protected
