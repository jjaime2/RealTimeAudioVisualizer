��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊F{���PK�R:�ϐui��3z
3�Sg��ý��^P�V�f��^q��9	�a#G���XͼC[ɘ;%�ԗ�V��-��^]�[f����WF1��-�uU�>:�9ݹ]�� ,s<}��|�cN� �r0�*]�SH���[��_Zg-��V�d��>���v�B�|���!�^���~B�1>�CD�-z����aS�^�r9Noq΍+ř�X�(�_�N@nS"��5��pxd�-/�Ng�������ڷ�dm�F�9�I�O����kc�hO@[�?!ѩqԖ�>*��+�MD"��xQ�(���1YmTu$f���$ׇ���O�����J��`�d~��M���#p�ʆ'K��ov��;�]�5	]J�W&�\7R��z�>��)�� Qp��M �/��T�H:�Qο���VǤ���r�(����jV�R���q�s/���ab��&����j6~1o6Ёۣ+*�`���	j�0⚃W���%���FJ��d>=�h�]P7Px��^\�A]/�[o����U���"�qh�e��ͩ�c�»��ܽ�V�U�������+�"�	�������޾i'!�{�*�~2a2� 
�bkˋmX��"��:�9`5��౞\	�4ZM�G����5IT�Giv�&��V㴠E@{�ʝ�Wm���]��F��,-�M�6~����JG�%��y�_`֋$�T�m��<�����P��r��r}R6���<{uJ`s�d��G�q�U�Et�dO�)� 9���hڎ���5O隡��5PY��\q(i�	j��D�/_X�|]��M!$w`�O��8Vެ��#QK�2����_�e��r�Mh�@����}H]CE�Y,xa�<�5��HD���^��3��`�Ί��5� �B�bV��b�����d��#����n`�.(&�HQ���S��;M@.�;Ӌ���4/7f�.�_�­��{�߮�_���5I���� #]��	J�i�����=^zt�ht���K���h�:�tg�p~Ӟ��޻-�a&�Hhu����ʆ����N��H��;p���x�Tnsmf'���� 6}g�t���m/���f��z��Ep�����)b���q4��V;�-?p^wK.��U�:0���^��� �]ƽ�.�;}���~���h�v[v��`�2���z�2U��G�i�3���V����y<ܤ��͸�O��y��%3#Y�g�o��uwf�TP�3_�3(��"���!�ʓ@8����c̟�p�$R�g�<����'����G��f[Y��X�|��g��	�ӏ�㢗h��i��: 6�-x�������J�ŀS���A8F!̟�j���#y	3Wǟ�C9�ϲ�m��yD�]�83U�e>h]>bV^�v�_�Ȯ�E�e��%=Sc�va�J�g�1A;���{�j��#���uk�-����\�.'��У�[��)���T�Vf#������-B��e,D4r��餧�v
2���u����c��Wy鱄��^�A�4���%��BR�Q ���^���*Vͤ.��m愇ޒ��(O���1=�׃*1��G����j�x����jG��G�C���+�}��� �ZA
y=�w���հ�a�����85Ieĸ��8��j�F�T��#���'BtnUYqǟS����c�T�M<C�1O���a�0���ّ/����[Q�rBLZ��_�ފ�G`zH=�h��(��|F)�p���M79c����<�1oG��n1"I�ۥǨ�=n�=����-��D�ʠn��֧�,ݧ��/^S|�e&e��)iE���
�˹�`�U0��=��K���2Wd6¹�� �.K��Իb!��K1L�J���"�G�=/��#N[sh �)��=h[��Ѕl�DR�V�{�(����z����R�_�q�<f�F��c���a�PnJ�v=��=�B[����VBQ,J�Xm�f��𝩳���<�j�,�[�τyɯ�FGs�|L�����Q�����n(L�*�`�?�:^W��_uYd�큤x��zb~��1Pu��p��`A����H��M�I�����*�'��S��<���x���K0Dg����ZC=���0-z�;����W��Zɤ�� �l'�4'�����P�Si�?�GZ��͈gn�+�`H'�gtE� �6��Ԛ���Sz����XAQ��a���:��|���av{ߌ�	#�3�!�l���
d���ިڻ����|�kB�>�C���"�6��+@|�϶UU�Ԟ�����1��7�� �|�Pj�^t8v���V 
�ew�����)uD���vd:ؑ$AN%+��Vz�3�=̼��!A	#����%߱��/n~�b�B��؍n�k�R5t�Z���-!|�O	s�/ +�W&Яd;V����yy��w΅�b���W)%Z�P��ؓk�.h#�Ƀ�F%ah��չ17|�j�I��d5N�t��Q�X���;�F�]6�����+R:���#%�'J~=���H[�J��+?��ǰb{���z����~���^��Q_��A�'%�p�~+ҋRz�{+JLظ|Fo�sb��c8s��r�P��4��Yx�>�X�<�R�J�E����B*s �	��L���K�ڶjw�ǧA�-�@����EBy���v�	嗝�R�Vb�����E�',��\j_�/! y�TEn��w[ ���� 3�q�W[��������^V�ķE�sf9a ��O�Ur4�=7#��g���m���R7�e4d��4W�#z#�YW�Րp���]l�Q���5:��O�����Y*.��Q
���l�'���'NYsj*�M�~�E4�U��� M2�*��8���nGzQ����۽\�u3r�9��Up�������L?BX8�1�uVGd����`�Kmb��r\�1}\�M�KwX6m��[����U�+�����W,Q�kdDpn�*�-�MḪa$*�ߢH��)�V�Q��/���o֘�A���(����A�n���eoZu�V��Գ9�伇������sV��b��펂�k1��;��Z'ۄO<��x,����/��w-�Qx$��t����ۡY��Z��D�t���$�h���
X8\�ݚ��T���gfg������RC;6�ܙY�&��ʨ�mLf/��2�m�2n� se{���v�a;�P�Y�w0&@�����i��MA{&c�i�M��o��DR4ls
Dz�^N]-�f}N���=W<��V����U	��/������M�
r^Z�����Dm�]t(U3&1��ֈt���Lˊyu�72+��<��I���^�:1��7lp8�0��i8�K;^� ��4�Y�eh�ny0���