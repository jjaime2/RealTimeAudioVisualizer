-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PqVhFdnviRDdKbwMTOUqNTp7aaMaA8RQV0YhH8/FN2htod7DUWYFo3A0cn5AKL5COs0IeuLWTBvW
4PGZDIKhSk1H526hBpqJOBxSIuw71uWQNqhUw9iLUygr1lgkU2/AzuhtAaEvnjH6t7/v06oPbOEU
T9uBTGyNchBjYB0Ov21IxdmMC+PD69PFiyaQt5lzC8aiXMxt0o0/wpYE0sLbMSQjzYWiwEjKml2p
JHcNjBMflmEajYLsB3q5qr3Jm3DksNEnJeQPJKLd94XPoC20KehpwvBNqfMLjQf6DdfzkXov3msw
DCk/jC8INsgXwRFcDz0y9IzSjPfd5z+L0OAOBQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 43024)
`protect data_block
Sgx4u4V9R/Q35JOJcNaarFsw4rcmNCkKKRLuXly96O208zmqM/+CG2l7bG1r4dh2hJB8wx9kG1+s
iDfy4DWG7DXIXaaMbUVM/kAjysT/BlamAfGCl2e3uOSFrl2IRZTnms+wmf2kgHnru1Nbtm35t1Ox
O9WDRwkqYbEs8PLj0Q/HTKxaESODKC/LiktM9UGqL07IAuWSnZLgvNvQC9AeFgynoHcq+4OqqIv4
wnr8Jj/iz1yaAv9H9LRkzrmdzGU0VUgob9+dZm3meh8qP24BOOSnVbFSOViSLHrUIe4eFQMut1f5
9CMUr2gBAPMbFesbdmh1TFLXOqwjWloz+UTN/Q8apDKDayqpW/o+PM4HT2aBS+c3inRxXx5Cl4j3
t/coLM0zUVeevX0BN6LGdB15eElKUkazyTbycgpJKjFSSJSXlrt3vR23mXZd6W6dDqFDpjdsbbdw
zHZehi+MNTw8iUT/ibZQLzcWfts3FPXlK4WNsfllz5thE364JFDF0SiLnoOUwv1p6+9nkMo5roYL
OjsH+gNdTc+xFkTks9mg6izTZqs/Zs1FT5+QipEuQSPAFVbGektEpb8kIWK8s5gA6Er3iHbx9eG3
fD5SfIRMdLlCCmjowFiU8T5cxWhkisweiA+CmrhjdkqxvYi9o3NEe6/y/L/vycK/WEeybGzP3bkM
B2VUjY2c9OMaUq7YPp0lnCoBB1XZuBbhc2mxKHkFGvBPL1AwliZ4x98xeL+6t0JF4ufXoGyAIiZx
qETFSy/OjfbsSOCP5gk9s5KaYBmtEKzMwxEZTX6TyJ5ZwMCU3mOt4IFytDt2mC3NlfiCe0czdO97
MRdPc6bBbCVbhFOqB35GveuBiP7PfHvnmq9nhtKfhvCMnTFEjzYovdbGvMoDEXyWn/DL8xFOLjJB
QbGZseV/eNV6CDeMHNtu+kdJZuEL7fP2LYHpUowcVhXKX5TzQgK+FRXqIeQgoG+cntvSQu9b2Iq+
qKt935hhFpSnRCe1NpT5pUninEZCfuFWQbbFi5EbdGY7o8Sccqllg4u/QUgxFsAFSL+af7NTgllp
LGHA/Yw3o5hd/uAItNYcUKNeDcwnJm3fYJNSj9SQrIQVZLhOyCFJz/sUPLSlsIujAc8ONPrv/SBZ
BNzIzPzyaTC4JKC1pbM7CmjR7dJmxVfr8uCyhpxJ8/p38mOnHEgO3Ys7Sz9E10jZk6WQv4Vn73cZ
+xE0+NMdAYPop3kjK68K/tYrPG/IqN68E6zn6+f3ssZMUB3YFQX65EYDsYNLnS71hcVIgT2eEieF
mOEQCtIiVFYymfAIRLzPOLy8nn2K3+cZWq1SOSjukFaGsWPIflaz+2IPM5eUh8GujfZX0OM0MtEh
5fGEfwmaoZs5efnsut9AJBztXOlvUSizdRbQIPPf1KSTg0kDqQzwtee00RTegAo0MQITWH8cMvor
J3iN5lJTo7tIEq+iyx2QN+GPFxofNxt88o48fpsYW+ROJFjDOevNVivAmriJiXNCfsttxLdOMpbq
IfmP18Lpjvr+RA7IiOLT/x2f4zS+wcYUAJ4NtYVKpGSplnsm7dxZtJ9Y2k2Yqn+qrYdRm/VBQ6mE
nzFfZwHpm5xqo/qhDKrDFFbvGkaINQKeI77xiVL3mt0kDhOptP7bzIHq9PzncUnWtVU8HMmvZC0U
X3fWhrDWVqAiiAgFhGD+lt45nI8ZAnqWMxwzTf46PlhS1kXlTq190MYz0wgPjl7Hh/8/pF6gv6Jz
kU6wfQIidAXa36Fw4q2ATCMwZP+Xz/kNjV4tjsqLuajTPMv8F8ykU7qjJ3HGaUAeNpi8CJJBCAAL
gHQq2K4UWv74uPqTjP20IDPXp3PFr1KFSQBr0XbRsEuheP5VGfcPL2oKRzBolbz6ZS4shaVBxayt
tqFvM5k7U+EfE6N1eOqszXGDAXfXwkicHut/9+quNJc2JM7uKKd9Btwk/eTdSnx1uSxgO6RywBKH
E1IXKnC86U5IuGqlQt//bNWPMS3eJe36oQu2Sui4tE0WL5op0h3MQerzwNnE9KVlhwVE+HGoz/HP
CemKxCaIbtKCa8DrngXJrkBS63qHncb+Tg0pdl8K3+U7WtcHb3EVXa/KN2l5K276xhlmX7yB6m1f
0IzWmIQrY0XpmaFJxyyFVkoWxe6v4EukyKAUHsV1hlU9hd8RgHMOV5U3BPR9Mrjyw7pVSLv/2oCM
8FzbGrKS0Qy5rm4hI2MZs2xafgfIKkTwZcz11Zoq2cbvGDT7k87rHEYbMTMS7izdmALllvGw/ZQz
3uLCZ+i2BqC6HF6apNDvdsvCia6zLS43P0UO2lqpTLofoVSYJOaZhiLbTgxSXDhsLHU6qf8vOUOH
S7MbONv/QZW8MwX4Fs90sIEJ0mHNT4R30rdm8OeQvND6Plz52zYm0cIXiuFlcijY20Zhir4n2ZND
kxdt5DTPpyeCBXSZzHbX2rIL+5ILN4pCrWG2sH52O50mWtwnwuQSTaa2E8vz1T5FOCD9/gRF21qB
80CFy652/hNMndM5WaD/j/Lv0lG8teeOkfX99Qn9MwBL9mF2zF7mIsP0DxHxPSQL7riW55Qz+H4W
/HGbwfGWswwq6KVuy+ZurnKHv/rJhKscAY9dxIJc2FohRmNcvep93XbWPB7JEuXhowCOCquVOn7R
HYpTCMu+S9kPi+SgzExsvJd2M19v07RbZyecBy74TE/04qSrsOdLRYSXJDiB2IBPFEW68Te7L+7B
9bT3xM/ul/SHiwECWNe7dinnXAh3F0aR2q1vfv4QtKJWex3SngbJ0XmNXGcZ+NSq7Ct5EOlcZywj
Oa+5D4JjCASMfCsjuzUeVYn7CsPO2Eo0tWniKIC2JDYTCW0dHuQz4NkdUaeWCbRf1sECDUCytxFY
GtB+gYkauEerhuMZBqBeEGMBtIqNq6M2rC7F3Z2SHyt5Ru+K+sHoY4xy0e4ls/tG8IDsWM18InjA
9jQDerTOmIcJt+0xxK3DNb5GSfa4lyRUoIviTp8uZPo0K9RjHziU4MZZlUy0ApBZD9qhXh4Q0hUd
fMiOBfzqO5xQ2rKmM6y1pqrDXpWVDNDwTvD5SZHV8F1DRHLEpi0ohKA6x8xhulHZDQjmuLmiKCpe
FQ3LBX0n4SjvJ+XD+HyJ7JAYnvU3GV86qQyTaJ7Oi60XgkXJNGWKn7TqdWbmV8sb5hrDBaPgFvTp
IHvApdxxfe5kxIGS3KS0dmLTHX+qgHYDqmyXvdsldJ+YlHDAD4v5AdeiwDajaFFyeFvMnRaKopCk
aNvXYKgC9tyQfHotSe1rjxvB/ntjCvDPaWDcNUWr6/A2xPW5GiS5hngybLITv0He6CGp3naOo7LJ
BLE228DzDADNLjszh6tEP2fOe9K/iYsIQ5J2o+/ZYrFpLV8PMK6tLBBhMhHVlS5GkzN4222Ot8l7
xmPZsIP+e4qtLiX9w4+iv5DaYfUOz0jaI0dzDCBx+cE8WCAQymL2VyvFbWboG5VvF2a96FYyfTfT
d8a2k1HOfEfNzn6MA4wJxNI//jqpVL8vc34vk1liKMNiMvsH11Ru7epa/JgckbOlcLuCKKKGe3kh
NgNnlk2/joIL8LeiSm3snBUqyQOsHPnZUZfnTgp9zrQIky5fX1qPT8taWsHwPqi6Y06T1anYomtT
mXdgwLNsyqKWQajcWsF22NXsVJNfbH69sl0P4T/bILPe/EzxqNrirFnVCCwXf1j9bHWsMQWJKCdw
geS6GAobkzRJFoNufq17rTdElPOVvL+qiX/wDfYXN+bJbTJp2v8Pyc+H1yqGLwdD4rwlrREiGKtv
bp3tN/lm7fc5MdaisR9HANhVyGon/XrFnOtHQ2g/G5qkHmHjPLJ8NBrwmelqqZkBNd6ogymXUqFd
X7jcEo40woWUr/HTv9dkuFlXbttb9BTQ2mqdIyulkSeIL8vrOQet66KobMnPQzY8CHwDnhEza5rM
M4tuF4KKTzGx7Hr2Dfq7RX9pXHayjGFHq2MqpKX2VbVw2CP9Kzw7Qa0rP9MrilbVimAH1/FmrjRB
bcvCCyACilgBWWwH9Wz6IJW0bs8tY/VO06HPp9/dOvSb8jgMyQBT5sLIQJ+E0n1A/NCQ5m+TXI/I
OnxvAcohZcNLy001YGhP/IYleIWMaY5IWeqnR2tpYTYBq//6jgZj0Rja3+5Tto5n+fZoTOoz7vsp
F14sXB0FEDsTmq2ZtVPlkj/vY6MyyFoKViAN/buEAt6Pw9Z49VJ/ViJzG69NtATXxgRwyFJtvYhK
e2/d1/8SXLcWqiSQvpEzMhNRvhDuruvoI4VeCLt56x2JjxnWXnHotZ5HT/93nX0zhIst6ybZqg9J
TMD+5PeMaDJKLhb+NQ5JJnMVouxd03z9cgRzgMHNcu69Pz4X3jVxygdqLTeFld+JulPfxqQvxXq1
eFPpvRvSRe82ka3z1RKq2kYCuf5RMgiiioYmfenlZOA4UslNRNyTsvWFrGOy0gI5KWTTwU6RS9e/
JhQXsU6FF0ZwDQRthzvBxC8Ra1o5GcMNY2ziUK12tpYCfEvb1hlnKwDdfXqGg5t8UnGn7vH+UkDD
GDnJewfeoaayfQz3bqThPD/aVHJDR/85tR8ZVuFWnlZTbd4qjw/Gome+ieyQpCTn/2UtKQP64LZw
5NauLTVAl1AMtLGSCxiaoliSHXKNua6wvOnOD++v/UOclTClIKhxb8hEgj4oJFFb9W+bbMZak3rA
NRTLoc0ZtH13yiUA7lUrosRnKmwJvujtCsM3UdIf48/pJBdKucxsy5JskflBwE+QmjQBehom86X+
bgc195+CzXP9/6sKJfGS5v6ZPChPHgcaV3ftH+lhK1lgdqnYTzC0FrUrhEtbkoF7SU+qKvrNC5wy
c+dzObAcxD1ZwU8+Cqh7XwSfPwH74u2RXK+GDQYQWsm7COuqz3Iw1lCyZAm6M9Rg3nNoYoiTcMtv
HxJhAfUkTKVsfH8ujNCLNDSpM+ka00K8kCvWKwywk9I3BqxeElMaTUCNLnrjW1bLyMA8ba48C83J
ZdDy8tHntCyzQj/nJKVWuSxD+hOZuhc8rbtsarlCV7c44RTbBH8ti7EstycE8AqXpsFReN0TTpPj
LiYaOKHjQsNcEE+UIVdSuemr5dB7IUwn1D1TrEoqUUDthT5vzi2LDbLL5+yyr1OBlGnmZ7P+exIL
B7cqByBjULwtGW5ISRsnOxvJljpqYE7usUy7doGhbWd/OxFWK8AtnKQ8tzPRPDbEIMqPhpPTqUeN
H3y5KeQ0mYT/nU8qxtAA1NE8Zf4Z1gVEjimXh1k7++mcHoSPS2LeQxhPMR1f81CHfMd/zQy6MQ5b
eAY5AbDE40ZMmYq8ZrY9Skst6n/5APKl4uqRsSg3hzbtgem3awwbr/1RiQUKy+b8cqGAw1XEW3Jh
GDoYGAYxhgUrOAvycphZ5IgWicj88/Czfbg5QJPnhO1HuGK1Z75OrV1o8ToYqcYO14MbJS51CdYh
qMysjPod1yKHGOP3Pb/dlavMHwqk1H4PbZMXiMr8deTNmOVRKPcTWulvLTcgjMcbmW3qDZVVfd4x
RrGy+LK1f2JA/GWPdayeZU8qYBMXNqRvJDkMZesW7q7a+7edvM0qKRgvvsWyrJoFqN4ScJ44p8F+
fe5OIKQxtcqAOdo9RBZej6sY2lQd9Us+O1iprshXZWGG4lmewCgDwWoj2XRpTG8fawgGcYGUt9/Z
712z2RIfop5Rqc0iBLdyxdv4jCbRnEh2xIyspDqu5f0G8SHkvr/GfPmdiB3NaHI7Q0nsvwVHeHk1
Tg/TZ01CE5ubrUQPvPjLSAJgkXWsspasyMyzea1VP3XjxgnfrJIPEWthGdqOEdoRaea2VRkiN0UW
S30lCicf+fCYryTfKUqY2P+DV1wI9jOEm1BjV3QuvlVURZ5rfU+xQYaxMeE1nFzMOst7ePggGzY0
lihZMbh//LDuCLPa5OXZmWOotPv7QWuSPJEcskYbVQOLwfv/4pLI60dvG9sJySkVHL4BdaqmFBHJ
pLrlPn1BP6qrzNI86riJh1Yh2l+JPC9dcpI4gRilS9zeCCNzixmEPcwcJ6mCigqc9EYjKtAoJy2h
ZPYt0llXmG+1/iPAr8bFZNY13S8f6jfa+Kso6J2nBfPd+MvqkQehEpZK4ZdOuruw97gitYwUFqKt
qE8Voy1YQjn7/2vaRzZMgdzYjoj9h3vKLdLnRjpVqTCP4xrTJ+iaAETzMEYLFZqq9SEkvGQYQaY0
2A0gQFxl8ZPl/o0NRequPU5E7oZAFGbVLIS06IjN52MmkYbOSFwFIw6w63TBVkJLkps5sAfLXUNR
4rw8EBJadvgP4wRLuPZQVlETrHUeiBD7Ihqa42lIYGBeHyg/qZJkmjh2Ld02jEZY+vTKR00z4STI
KbOmIvXtGZHE3tIE32sFm2R7az3macyJ/ge+W95zFl0yGRuQ3tqOnwS/O8SMj0bYOFLamQRv7OtR
Vda+1kBBpxr2AEBnzrLQlFeyM4oAEYZ8CA7oOp7tq/njYBwoVXCgrCu0FKdeTR/v04ueaQsu9cll
IdozbtCiZDvYUWaLYxcGcJK7yxYd2gGQwAR3T7y1lzICZc49vWUWCxaQlQm2BbhmmlPqfv73rD1q
Ha02lMD5oOByz+fhlR9scXzqG0GJMn0uh0+elWfgK2XhkTLw2y+rWUYGxAJUptt2XUqtsYOyE98h
+s9SK6eYLjuMYB0dpQVueFmbQMfTtQyrXdY79A8okcCBwQjQX/RrJb4jBp1oRgO7jKbo6zEocEQM
5atStP9FA0xWHpy9wt92D9zYhOFUXQIZfKwiYiJuXSmUrFxlamTLTp2pyiSJvjsyDHPfEFOuToEU
ZgI0zQI76GWLMNEdRFGwyNyKBFxiMB1IhKWa0Kcwl0JNRrsX1eMyhUVL0V8JgDYPLe2IYntk46W8
jyiiLQ2PlpC2cOvUSTap0CrpmXDyyRBu2+uNXF5pvsm44UFsgaob4R4PWd80HS3xc8liLCnxgN5B
TpDY0884q8tagzUbSAr87SRiF83mv3Ma6liyjHN0IB2Svfk6q0eWfVO8PYaBG3ysIDT1JKZNs2Oy
HU4Sez6hYOouoesOMpGITR+gW0hthAPf+sHok3wzmYCq/QzLCxQ/tEjlWps5M/QMFLN4i456SW3F
GVnLPAgIhRVfobZmYSMidJJBJOBKYQcxez4s5dXayWvNFYuujYpEfrsWFZqMCRkFvKImIh5HrTK9
Ck7sLkQs6uwRgCIUo2RqabmOD3a1DaaNNf4YoDlnA8EB9MRXOWgWTgfclcbVDlD41boV4Z8i0cjf
cZQ6VFFtBIXqM27ADQbaY2ROfBBmrTVFKEHm33XLaPgYN3l1GnMATfuibIU9s3L2+qMI3gHe8w5g
qx/KasX7YjeBFDph5q1ujQjhJI20vZAuflwjwQns/m/ikohjDkxGw9h3HT/ECBh0tHNWxG7ztpC/
KgAMjRibTAkR6A/Aaj64IZXk8sAH6i9uyvPRFiRvbqdJEg0jYqUlcIvfuIvfD/uaaVrMmYXYF9rs
nZT4Ih8xXjAibzhmmUe0drDzAmfyZVxldLiKhCzG6BquWVcMLwYdTHuovPV431bAALEXz4Yk84dY
tGpN98LSz3RJyTd2uCUAaopBIYaUZdvvfo+ix3kKhBRqguDIH5rnHBlE3yEGWBzyr14DFl6nzDiv
LYlhQGy1p//cWhJqNmhASus9+LA5v0YgTK3tJ0BZnIcCtUIWTqhoeAm9Zt7c9dKBUv1Qu4+iwHc0
Y9zJe1k66EW/5DmI4EVPFMPF6/SeyonuzIi4ip095dBxPLQ27p6plKkGOvyMqcxTeoZFGSjdLmDo
6kwWetw1bQNVrz1IFzKRQfmm/WVECxg1UkAHGqpZQtKBR7rerynVdDRe68jhr8kNoFfsKjf4k1+v
NRSwJLUR16ZBBOBmq9l2TMho6MTVbZfh5GI8X6IVHcm7TBASR4t5ekxSWHv2lrKNmy75f7F3heYQ
fZt9xb+2QEBzvaImoRbRn5IPc9iKCRNJWau0mallW2chux6f9dpGn4jJcN8Qkee33F5nlk20tBlZ
K06J0kYENeVidOUBbtwHAn9SA7NUMlk4Xxf0mJbPTIj8enmo4T4UlvWRPHfJq9Oj0cdZPVBRcnj1
V4rYtP5+uyNXFbMPhLj/kQiJZ5pG3Nqmk0DkTOdtfGPl8RVziuoJkSFkHDzXj8e7PHHxt5uW16Ya
i7/jeJ08DaeNPPRiEeyvmZ13Fdz7XHkmo0YYEYp3cc4HeKSrKN7kV6JqHoxsbI42JkxddXPrJXGW
Pu5aAXCUN1B7q67E9tnF14qmjakne3UFGUSVETuIdTojDAjxmU4UVCRaJu7/bRNXE7FnPhdNOpja
nGf6NWDt6XTfDbAyJa0qXc+yZ2KcmpoPaSS2BmhnhgfxjwGvINOV98rshfmc+kpO9MSZGZrF2dGW
3noP8j0b7/6EMStIdjYWN56/BbmpBh9g/qsjfAQzP1hQu06QP8CkeDRfPIwB3NL0tdHdAPXvIQEf
rYTGVnGJqzZlctMjaku1PUklj9D2HynLfDs7J838i1yRt4QGnhNaS9YxBA7rFNsLyh3igsBcUGRN
OCMNANczPLeaceyHwa5YUjdLX5POLdftVGKjFMeerE2f5iTcf6ywDCNsqbFhIjqByPa7+8sH0k2g
wDmRQMjoBGFLwPqXHdP1Zqnwwxt4fs69IDfG4SkvH6TAUJtWb/OuDgq8dPmHBvoJG2d7eb9BLzXe
TAW5lWsfNh2TN4bLa9Xp3PjLUvEHrDvfvyUQ1+LHjmbAvMUH+zzm6FWyFHLaBQWACIVtB9mHY/LF
V4Q6wpkaLm0moasKh5QhvwqerXdwkm8jRMi+qeC3esekAFN0jHWX55Y6SPHscQGa/HKo/ns/PCS5
pmO9esaNJJml/+8MAFttB/EMXiUxjxv+c6WOKoSGnc547oLF0q0Kde7FunIlLqxs2xUCXhdcnLG/
n4k5182wgNFIJvyaRWcq6b68doi0BE4jV+FzoBnnLKS6YSPJHQto8EG/hIEI7GMFsLxSqn3W1DUy
6yBDvtY2YX/eyQujRNQ1dPbWfDp5GxgnHh/lH9pi0AA5D6YPUDU+KKQ6ZW0nDUf7DgIUXfBB/n+i
sNOBNLXZUJFiCwi2oJthzoFoP4QyKJVZrBAXyfM1rSI/hKGbAO8HbUBvkywcuwJxqeglDxEcg2Ka
qtn3vejxEfQI1+j4/FuCdsrWNl/Irtp6MokW1fsaop5EntFFzwkVFM9MgiSdLLckeD/2oY+jDGnU
sLX4KNjPWb8Trf8K/BYpaMQZrdllb/xfoCp/IVj+WvUIgby37jX2QuXQ3mHs6IqW1/7ZqAtoJk2Z
qw7rIeU5kHRKlcncPBSmn6NuNSY3D2BL6U65FKQzyIFdzqhClhiO4KWt+171ifF0blKKhBKeN0yP
ZjT0Yrmp5SOH2nq2oJbK5QkszDlnnTZCOWmv1y48LnDPAlIaeieOzYfvVPmRoPho+ViCywvEi0cL
FZtDZOj9HJ4pClQhv+RESRvGFBWgTNJkaxzzfqO8rhpgASfB/0jwl8g/ZqD6D9iksfA/y8r5rRuJ
oBSOeTurqD48C6Tnm06nlD8O7cg0a6H7ub2HLkVvdzJtw0oZXd7/tpwF4HE9da+Qe89RpF6vl7Kq
GLVATNjYgD4zP7LoVGA34lhELGEhCUb6MMJBAYFLh7hSKGwm9mcfKmTz1zS8ssm2730wrH3m7+uT
l0DxUxWlJJXNh7M6Ilnsw3Zc0quxQS+rLN2uSIzSz1TBCg7i8Wj0GyHP7cf4nyZhe3sO3IQElOFh
CslMcuSv9h0Jqi3def3GAZOpltPps3gmyfDiMspRT9QDTc5TJ5aMDO8alX8r7C90yvhn3oH/xuBm
nIK9UweHUFlw70xj0eJH3yPcPhcvy6Xgnec+DaJeV61zX6okVuZUqODVsa8M43SRsMXi4w86qRbu
oknnUTPGRwPFqOlHySkO3gtnQutLu5a6I7okLZ6bBDNCmla7lZPPIh0dWJpNNM97QYiT+QLRfahz
1oPo+/Jicp4VBwi11oQiOUHVVu4Gh6ZvnOxQeQFrA+u9NOu2pVMExfM8EeiIUdX2MGMadDJzqXwZ
uGTYEeL7BxQtPDSej4irudKvnCs2AuZclXaoqp8g2kqldHSloOPRxhNx8E+Qphnh1ugk03v07F7K
weH6AEMByG0gnyfCpn684hAtXTpnhVEY+v6/sbGbULJWn2TXjgaN3zUkUdNLot7Z6ddgTGoil2jo
cqxAjsRztTtnIe5j+3Fo5PoTZnf9GrNVBLBM/OQbhH2bNiczKtWBdlsrzJWO33yu1sQdK9N4KrDZ
SCt4XraCSg544X45y1wn9/6vV2VtoF8NDQwAjqtvx2q/Gl4KQi6EkIkIc4m6RyAw/99UYpXfD5mZ
9YOXV2W0s5Dw/MEqw3vesw89yZhjTMt1vDzdDKqY3q1iYRNdIALPvj8hRoEMEt50JhVg+kKRT/d1
er3Zdx2bz4Ay9K60D6edJhpeTSIghxsYBI+FkITM0yYpk/punSoZj8UpjD6oWahRIRNVcGaV4Wa3
a3EzhUlTbz1VEu9E2fqic1iW/Vsswl/yiM8zRqeU3MdwFppzL3FO7dS994IGueq0b3eukpVMV3UF
1+hbIwSnVqOc14HZByCIEylClzq4cyPD0FMm8C95xUQkJnblTakaWco8aBXuEMsY4MLicoamQGpj
XMIOLAHSJ8aIbqeqqj07p2NQq4WezfS1vgm8XscMfCxArXRNFuzmtPO6WDcVrvONnBwCenim07KL
GF4lJ2POe5RJsU8OGaqTYY7uBDqKmvz35PmvK3fEJHpasVQ/UjsGtsDmKNkN2+lCy4eht75ifVL7
LdcLwZS2cd4b2DXNY/YszAE3/N/9xTrqivtGal+6W+5XG72zH4+TYHe/eLc+UA8aDS+dknBIGPBo
1V/HaMhPtbF6INRiDDNbnEYDKEawMDaIPzQ14mPMsCqzyiENez6zVPAeLj7k8HcjQYPHVSL9nrdd
szWvPprbkpErcgs8QiyR/a3SXpbYowfvhYtGoYPiy0LjyPj7qhBmRW9/W0dQuTi93Yuiw/wyzZ/J
e4eRwgwwqT64f4yONI1KApnRPpzyc7u65R1cHiQWk4ZeocMjzvsOISvZF0ivCYv5ToDv0ie1m+TP
rAiP5tX5FIhHTMH9lADFCaPvocVakbX4+Oo7lZSa3wAD6pTP4JxPDapHKDA75MneC73DjcC+oOWL
su5u39m7ix9RxVSEhKxTFPqjjkeI0OL6D60d+a9NCXb98+PJ5OM1+KBdnaWTNahW3wQMS3GL9P1J
qEwr0B+ZPJiI+AwkuR/2rfaWC7sPqS8pI9xtmhkmJ75kuc88uonNh6jJCVwFrgr9MZKw8/tIwzjP
Je1NOg/lyUuaG7sB8+EIviWU0sWfqoUHRGL/zFL8s8WsniPMAMyMsA5D/BTxVTcoUHJ4g/VhMVuE
Ss6Y2qcL0Pvg6RbZafzS9OuqHLoqCtz24Q9vNGLD7Yw9QVlT1nKlSDi2mdvVo73JgdlYVnNSrREL
/XJ0kM+LkHgPAv0TjyDky/s+PSxoK8i2tU6ZYhhNNlLZY3E3CBiW7aj5AMl45w+wFV+7mPpMmGns
qMh9BBGC2454mJRMZjrHBgT4NHWtO7THu5Wfw6NRIPsNNtX0AcDU7N9A9MUwF4VawNemskyMDh1C
ASvwFKQv0p3VOWHQ+OywOaH42hXi/qtCufy8Uc1LYLiBA1wL0K+pZaRTUITK/PNFYBeueBnccanj
5MYrG4mo/MnhBTJll3wUHEufWzLeOdXInW2q3VeohhjZKtJELmur4z9W+ZeN3Z6E26pGgwdMWAW1
4J/ZiUQeL063OMLQg+MvFiciS4wWMKbEdKuVu6kJbxdW6Q2GpvFIVmGlA8qNmHWfmkKRyw+jq9bl
78EAIL47ocdZ5tcwCXKEMtTig7RtJGvSigkAgKfd9eVKougYOu770Fdj4qy6JtdW9LY817MbOHSt
SF82ShwK2dAtLOIO7geLaYe5IGgPVTzbAhyQnEMn+sJG43bXhjVwkBdRc/tjioZVXskjL7A0Pv0x
mwZs/p3b/TDUBaSy5Rarq57aEh7FHwE9kzMyZR++vzgAN2xFk3UFn7x/zHQVQvLpn7GczLoN6g5t
vlnTDGiUWiUT/FFfMyauyH8JSTYw76tQjXeZmVvxqdasN9tHOtrrb2VXaORcK5LPoc45hQyMpoQO
NWfUfQfUDunVlrVZ16OXo9oL5YN71OUJJ++SAvhjRWt24Mx8QQZDBn6JEmLbCWboPHm0HT8MjmB3
2AhrpSe+2NkI8hJ+iF8W6lwG27gT3oqWT52CV2JQ7F/g6g3ZtgaPwQOSEa9Bc4EojsKgXbFIqoGf
AWLaOqBfdjIjQSVVCmSYipOd8/F8eQ0WeX9LFQdFDJzUJ0rw4nuOnwjxTaDmr8RQraBnQsQY8MnD
oHb8FsTtoRZaQV0Ew0oW8F/ZfwcPntVhFHDXL2VNlEpMwWvJNBMEh8/VeS8n+/lyZPwND3c28p5e
jf4pb3zkNb92qCI4Lwr1sDXE1Ox6NAsS1g7YZ4qvRkSt/zXTRemk19TYZBN5G9f1sjS9SkAYSDbP
WTu3m7+uMFe0UElh/MA5X/HbjFPDwXVptn22fb2wWkRqJaUJjLLuxyeJV0z/6uTlYQzTO7VfUi2w
rNg7nrEb+m/UTqGmqZEjlfaAdqH0KKVDxI8il5GMX5Pn6qqupDXGj5c0p1tZj64E5OECw6nHc4fr
QVWylA5mW0CjbinyBYkoP/x31PFiGvEO/kKxtbSXh8tUn3kamOFPdqIMSmvsgOqDLhnVgAUHZZhU
PC0BqoY5ZebWxZW5dnfn6G5CHIndxPYuAWDQJerOrWo1z674iVqfaA0qBgZuwgMNHe6/EBOymHBr
77COAysDUyGyF3TKJkKDHO2rkMzGFXzwGDQgvUptzgf9ZvJ+Qsj6Bvh372bxSxYbMwVdFxB3gJ/v
O0JvXCpXteTFizvomIluISBWt8gap16nOb9oUJ+go+Nm863rZWUfU+GqI6UjKYHQyUHQydjM+qGG
SUrKzGRVzy2X+uwOiF37GKP1+6C4a965LgNK+Hi5LOAuCrTcsvwFLBvYI0+SrYX95HKkpnBbH1SM
C9+KGFfKIV5CMpteE/UAutguGQvhuEYlJ+BNTxb+iYBWXMWDaXqnpk1Jix3CciT2lK6FLRDUodOE
OtEu6NKc71ylm3XMJWPGi3o8msbSC4ul3eBBXYdAifT8TJM/sH1DSAAxxTlIHpfOQREtRigtxtVR
UJi/DA/mExHZjHeijjSyjAg1ahmg6RpSsKrhFQeKwdJe/6CxrOgwAITXENtCN3ofyvZZuOreEJDi
PyqI/MYS3UqGbILbAuuguzTEwQ1CVdTcsnegl0dcGlNf/oP+IjI2MjZ5i3MY6aByh6/x7dsR8ASw
LiTKq01w6kpoLsBysrPaOJWRWr7vqj8pl+AfsxE/uyd3Tp4GE4Betp2AeVb10sAizNUzECc8NlM7
Eb47/cIRysYOz8IANOk0bc4jIgVw2vZVsh0tHP03GN8WJYAprlYc+g/U155lk0Ch26jWEquDhKbl
5/UAl+Vw/IZY113HocrfI1mNaCKyc8oGfi/6kNAIrQshRxPoD/G17fgF2gJiLVRxMZvTfbLmPy+q
+QHmh4MgtLG9LEa4+F/7LVp9b9IImjhQmLRpFN1oo/9FYJDUPO4SMSgfsKFdZK/X4JG4uF15RwU3
7oxd1gpdcYd0Bzywj3jljnebvkX10SC89RmEFuv0K8VRYOiVxV0/iu9kigC0t4MhmKWv3CT5jBrl
GItvu4vbMiX+TtSzzKHz8IapgwUF4ohcON5EFhPwAP474Lh+gvVOhuOYpK+1xk1qpcfMQJBVki/2
FZZdapq/s8Y5lzQ/xnZSYRzx3U+ngihqsj/0KJ4xwGVE+OydPJFPXCQT77KeOWLvj6ncWlnAGx3f
FtTzjXfsxyJDwNdKXX1yoWyarqtWCWWVsHIRFfs4k7nCzBFUF/JR1/1EDsnHzzdhy6nxr4UL0bSN
XJYFWlRKuskocK7CqxdHP5+jdip9vnwC13EyXBLWxUwtsL0oPNu/AkuaEpPHx2Iq3Y1k0AfCw4f0
5cV/xWFq//fBNg2EYicZ6A3WabjNHrBrP8zqyMGU8szGBvw2x3N6DXmSnUUYVkFvCtrOd8B7ujfc
opr27Nu/i4LKKHKJY3G95JfqXVuIrWLXdxEAqSqweUZumw0Qe2E8P3ziJpngKh4GxiRALBokw7Dy
2ozHmiQnNwlOXpMiEeTRwRpzHJ6DB0h1i4EdB4EIn9aVw/IfklVOOHLspbwKYX7gbDBF4vGlgX5Z
nrTtnYsrZFA4JaQ8ZOjc5LbQNOWTPUIcpMV8JHcxdtswOWHvE9/gnvfp4aHwO4tLX2DEedrEJWzj
OV0ck4A7HD3hnXVIYRREouBVvOmMbf2Rpvrv660vZ3z2HpJ6eIIUzHYycxiA2pKzSiIhieHzNkFL
6pDWQz+2ILbgPsV3AjyeIrIjbMNpFckJxyflNB+cdwSEWBjiz+hDvlmr6rUqPw6bKU57e4p79Fi9
3T31nUrdyqWV/lp7rlgBNpQvFs3JDdztl4egYyy2GhXlYslf02dIN4Almw23cc/gJbUd1Z4C6TpQ
LmUjBwA2gBTZzcwjiYZCJHu+SPTOUaFntCRgi9Y5SGEn22RjG0KXHs0itlkakB4sGB8Zs76tke2c
QacvlK8GC1KF+0O4QRJNvR5SqAuvbZy39oLBOLMx3PSjZMjyok7u/XgKVq40gQnGmFDzVQBKZEkO
6hGRvL8k476dc9wokxtRELRaS54tXKF1anPvKYw6bO463Wk7ZYfyRawqkCun0YLxuX3bJGcj8nZ+
N30YL8pinEZkRKSnR6cf3v45uR4WgFXdCV808fYNX/BW0j2NGDBmkFD7lVprFVeNFC1DamqOX9Wy
5cmUG5La8U3KfZwjkdXnTw8RgAeUmIZQ9/cVaEsrVORKLeOGmdp3eUYL2TWBpaGOc8RFXDyxN+t0
CBgkGDWdCIsRh4J1hQ0/uJ64WCeXDhreQb5WAP0hUn/uRzzivQTH3xBSSsCbWqWbav/cY6lIpnG4
Q+zzJ09gdUbGr0OSRQDWMXhCeJB9vWhcjKH02Wyf3XkKoMIZ4I8z6mvHZc01sHN1CjSeoiGRsUaD
3ttbHZzwIJ1CQ0SUz5k1jDwoX27cPSEq8j5ckOyR/Xbx37qnEmuOq7BjYOgOxTv0N9Qy4bY/SjL8
tCPgtYW9gxWMzwg2ppiLOOZ8h82jq53HHgGU6XVyIzigKxXQpN2i+mzyjVe7gFjGvpgmIHH2XVuF
04nrwfWbrRxCzwVQ/7uvNDYPQmuDEA4IOD2DYklKmMVPrEPf7z85ePLYj3wmYMgX9cDWALjZzurb
mwmDJUxvT3kZ3L1Fg8UMI8rAbD9CeFoL8Ikhq8H6MIKVuwcbkpEOSNxVtuMq1L3UkF/4svicflrQ
k2V0eahozxyPoWQjBZyvAKFhgdTvQNW+rvvlZzIkALHkNX9XDQelAEFvEt3jfekxt9/KLm6yXdo1
0GlVz0NE/dXCAa32BOvjLCJOb3LwLj7aNNYLUBKoAlYcsymBvz/R+vQDuMyURrh6KIBBacv0K4RD
/LtXeEE7JAlq/P7q9IpA9b4UnxcKy9XYZ950egyrEinWUM18IDUSVJj4hCAbIR4ovlBOyiFcDQ5M
uLxGrASvdOCrYQ251Q6+SQ6Olcw/5fh2ZSbcsbeNpfynvReVeOziicVH0VreFtRCSvQj92YxgtXM
skFEv8Xx6S3ZFiOtADT3XjGhDqBnK7YcQp68Fx2nrn2feawoIQMlpXT34114ZTmTDPYDlMwSfK3u
dD/YtIvN856pprIwHxH+dSwANP6d9T4ucSfklfglQT8ALOK6oWeOydmTPsCP34T2MykDvYim2HJB
TlAuPHL2kI2E6w4loO6nskchz6zxBebE36SowXsoTWZzgf1WDe1NpDC7wvicm9X/XAQohXzHFZWt
fy4QEEaweEfYZukjWx1JdkkjO9PwYj1C9ApOMk/ZBVpJr1+qSBiJLduXxT1XrGa9trF2wmOvG2n9
ayoHmKWdvLNAv3mEozPCnrC6JsR3YKULcEhxjr2IfER4022q1H4FYkXn1wgDkV3XF7+oZ5ZCbgig
UcAOCmu5YcFjZVTI87qwS4DaRZx7G466jtEzd8zRE6GSr+hR3NuOzJHxzQs6094B+SviYmEWl/vR
0CyDNoeZ41XY1lENNfaDQhf5gr+646pmzxKnmT69c0ma2YuJ8lYqe6cZkQ0vyHK/RrO03Cd+k9O8
C6+koJ1St8Uhcqnto0P8X3k51mBGzSv6JvdxSzGxVafQuGTrt1cP0f1UqPWaRiDLVLnwkHwqYJj9
kRklOVDpiWb31HQHtJynK9pxRccI8cMJahUqcVRp4ToIO3RvrxlFalxBBeEb8TlUAgOJfDmUSA7/
bSt2cAStQzpwBZVxKoURPBOEYoTSmHZkiLrxcGepWgAkl1AlwcVEOctfk66g4bPZddVv5/efOt8i
79b4JEDEncINWfmfkTMo8FQA75yuZwQZWtGAHsFSkxDYZnM0FQLN9sBl8fSi28xWIu//SNOdzuKG
PSgltbBPbM9qTCoUXeOYOkJ8lvT0UoVI71UbXmevUuUTIkwlok6GH+MLw18ym4d4vofl5YpH577q
ZX08W0RoCR4Dtpu7YptOJtsYVJ3tUnnbvvp41zeTZ5d3R4ub8z+V//udHVBqssqa7UKPyfBvPaS5
36Wh0/bGmweK1sLGCaZc91PQUt3ihTvFjLR08w5CpPejYL6Wk2J067TU5d9xgGQk+xu4k3cqiLF8
LB6lS0Vjto34EVJJ24INK6WSscQzaywm2Txh6vs5QSvfi6qxVI1AMJ+7Kh+qcVBTK0CnymsO4e/G
doswZ+F/3HrRqAWsn2iaGmRUHyvahJhVcLjyrQzXfH0zofmSxDkGkkUfDtXEB9KpYeFD9tJCKK6+
XAp4O6no+LG7vwbBhAZAcvSOW+WMj8Zh7Gs5ft11+7s4H3c2qvxRci9KEICzlIUpVKpFZUKATWDJ
egbqXJOhLmAZqghtpZaEC5aTwJcSHD4io/mrCqaII/+V0ThNm59OMNIVR21Ys9BXBaMdhE+Q4YaJ
GXbaVRR3eTMlsdQ+GOFgGUHpxLIedTTZmMCbm9Gvs9NqZWhZjFb1Fm4ChUhCb1meOyWIZQZWXjfC
hqC03Iy6glkbVxCLQNCDegwPuV55gHx2UIIBJK9Ie6Rg0rVcAYPFXN4abcTgy/w+b6NCx0KLKMQ9
1U1siry7L66dfjBA+lc6MmxQS63kiLPlrw0vJYlxS2F0PipWIbliFytYvoBhpC0Fk2h+pc6/cmlk
w1KTl1szNRJInE2buf12AWwVanL4REYQOL3F1cnD6h3U/k3BBnSvR+WgQBRdKXRZlwHw4AhN/ygq
+yoCLX3BQIqDUDPudVxIhOVnB163+s81iCiyNze/BqR2ukW4ssnIUVlW6Rlgg4oULQuoyk5tlu5e
mBrCtnDcCRIJzfK/F950zaDrx7yblO4INOh5Ixbfr0Fm+fjwIuG17/afmgM7PHbkDAXi3PbxecnU
2EjmVtVVDDnR3nAXBWD4dTPRsvzkSlNg4gwmYYFjrZvGTyfRfB9vh8jrslpV/SuWnF5f4lQNmK8h
6I/Ie7ERx1hgGNyhUkPM2JrfHOoQ9LHzF7cQ7qPri3K34+bWW11bZbrRwLXw8WiXEptQdnoIj4Uw
ZE8AFZ7Wo0/icEXC5UtjASVVSfubxwKV1lDiUVyqv5F3k07SpHr5OPutYkXYQVo6z9FiT42AM5eN
OFqaYMXXKx8QySOEF3zZeq5eZ4eVZmi3FloztUbg0HEq8iOiDWzP6LNJ4SKbBWnN4+FW8fIzhFvx
KPFTcCGmAr27veNCyh5DqZHyE922IOPFbzm4vOHfXx7QRFDiYmKqmCM7kvxrazuP624XnSLrX2cT
MqgKmrV3J5T/RFXBWFlrq8mfPUG93TmfiZTQyjHaYHEeXdYT4qQrbD8e+8Ur6ZemezCY5tVd+GKh
a5N1Tzx0OZVA87563LlbQEf0GQnoKnDQUvx4SKcaRm9Dqid0UiK3Ylw5ONsUrV6bAwypRgpMpcUA
otK+ARPKKNiCNuzv1Q0vg0OUZTcivdpfE/HwWnUioG2wTBLuc+wmYLJLxh1L+Xx2vacLRP8jG/jU
S65z1sep4YkYEGPQ1Ajrypg8kaRNHaTT1ZMLKhB02nAEka5Vw7ZbPtPBPPR4LuljghQgXzyvPuUh
Za8BVlSpkkOdm8haywtsN7ejBmsutMHhC5p7fGktZrV5WxS0MfBhbIhFR8n0GRdxhu7m6EQeCmTV
pGsnDRI8V8geQLE+Xfr0U6wDeKJJnbVbNkOIEuYeDn2EkU+FU2dpTIiyBhNW0hVqi5iAtEe/KDOd
zcRHK3hgmbSC9gtgfP9pwSayx4hL+3LRbsJiZtGsgOsKDQgCMHxr7cjYFImzcVoh26p6bX6VyI+N
aK4cnT0qYT9ic6Ln080kO+6EQsBhNbptJQkSeIAfGqIcgLiOpQ9pPGnYAgCALDO8z9D8dq0wJEId
iIsLLzZO98g3Sx9dpKLcQNSHztzbJ0FKyp1Bw5qEnbognvWLToZwyDS8PYPvlx7YwKpg42dP50nA
oxE3tX/LL9gjVyn6PtH6k5Hw2QSdtR3igIvXJtg0/+p1uaWNt2WUhP+frl5hodLEO7J6wy2/Iwxc
KAMLNRT0TzirPvYGh+N3KX8LAoTMO0aTdY/U7k8FU3nZMI1WkuuhDuKofkWdrTyrUr7SczUAPADk
+mhDv3vjc02hjRLfAk0WZ6e/ylLPr4VpaPElhuRAYI6IWrBHt4tZ1XzaLUiH11EdKvCKLWYVzoge
qknfRUKyXg7y4FGy7PRpaJGXmXpr0AMp72EGcX0hyWQQble7W3lyjYimgrgQBJv7HciCdXHX4WEa
U5NRwev5vjy45fROBVhnZXDYbsUREVv9s6G+/cWEsu9RBOGqiBs7iUOwqr5jEHN9EfmhWa5mNg0w
KaZdgsCiOFxfyDm+zUP+Fz8LXZ6xBgZnd6cXEF2kkdxTFRFwrTY6h0Y3FUQj2xt4661tL8QjNfUM
eRbcxRqy8ENAS3Hg48dNY1hiE6JGX6YMFspbBIgPIbY/o9xQXjJpDx3Dy0ocSCoApD26q5g7+MtY
3dsXnmv9xothzWlD7ToITt3tuFcg2O0HHqLhi9p+KcEiCoGA0kcb3Gamo41PEkVK2ho1WqpcV064
xTfBJ5aD1yf2lKtyxC9P5Vlhlbwqo4XJN9XjmDRwCuTx+drBWosRpsMtiKXXInwEQvbLkJqL9gv9
eb5rHZyHtMpNOTkLYdZXX3uvgeuga0knCFEA2t9lmLdX4V0hA4z5i3FobPjEULOgDmNZIrIb02qA
YDqTr94pBPQaOls63lGCorIZxkFVYburDIZcGcIABYNkwUHJcpSXrbunyuvE+MD/iQmLihuV/sGh
5I3jDAp+63qimj45naulkDhX41McFl7mHtVUVOQtSBr4idC8heKNfS6jbY6cExMEtFhV7gOtrODc
c4hvm52I6BT2A5QIyWK9mfvrLwOrAZzqwDMw/GectLZaKHVp8UiP3avAs7P2t5TIgSlM8UlOINUz
Bo/DvX1RM5yTl9X+RsOpHWMuc1mwTG/bx8WePqK1xaa0VszcV8MoSfu+EZOoYK1djqr2WCGnUMoK
45ExEy8fyHJ4p3r0CcfAEN/0K1pWc0XnTUcgVlwDijCydLzaASeE7XObSrCO/LZdGKdCCKs/szw/
6ZhkTGNJJuL8uz1qWA8Z4lzqz9NENHjCAjyH4VAEtUIWWP1rhXOu2eJdflYCuU3MKssn2LG/cqpc
x33CL1sjewD85cBJjI2Y56ciEIjbZ6YRVTXFqqkO/Fvlf2u1+ge+bllkkwHd8gpzKllO6uwnV0/7
tRl6Om7/iKVwQO+Z2vgQsFwgIjToTO+f74X1ob5k6cvvKACEcevXaJRDn6RnvTu6n9LFJgzxBvwH
a9HVIXCY1mZAfCMIZ334JX/j8pBWWRQ/CS6I/V2hczJISnv9m8Cb71Ax82FUAgntaIXBhuvgj2mL
zOZ1VCuOJqEPMkAG1Avl+s8zo3an9E9gkF4qAwfkg5tyMvA/DOllnc2yd/3Hp2/J1SctoNL3wnkF
5ISOfY2Ta5qTA5JqnggvROxYj01vsEyU/+xJ+ddUusHo2iqpXku7ZYTp3HoC1O+JAQVj3JJP+pUN
+cayHTy02OBaiIdMFggOUMKLRvpz5VGQ0VbJ1JiLgTikcFasy2khI/j4aAGtCdq5DcaTXgiGsPYB
/5hR6qEjDQYST7LKvkV6yO4JZsErGerIspeC1b0h6c0BAi8meFesngdq9aF1VF7E9H8P/F4uOZpL
kOEOrfvb468k/y7mGVXNufiF/Pm2+q9rMHvceOmjDNf2kz7I3k1t9cKEvd5/NMWp5K17u2hdNeJ8
wuW++eO2hEgkLJ3mhhTF/ttaRXljKLH0hoq+Zz9k8OTMNRv2kj5y6/s5xVq+3T9ZsaWN5li81+C2
4EE5FkCpdB1+KfwWGDsafplZk0wxFes9Mpkk/oVY3BBGaPTPYS2ueL19pXpbyptLn0C+1Xvked39
yXgtU9quILyffMAaJDE0ir6+yXEckBtuz13aakl2VDwfpLEylcNCkHmWWkbhY2B3H2w7VoOZ1gsP
zaSua1obcaM3WEk0qvq/zKwKfo1oQgrk77NadcO2pC+tAo7ofqImKtIiwBFnoXwp9eWa1J4Vq53/
xysXoXoCmkhvQVRaSKpcvg4nG9JL5QQ3v3Nux6k4dUN6Np+8IhmfUZv71u2kRAwVPHnV1pWU9hw+
QAgExrxoVl1NUphAfWVXUxLnlZTz1Z2mj9XEX5LFHqnqjDXnnhOlZC9aJE6F/xphl2Iv6subRhRI
171qUROs2eMiqLwiS3uMjTCykF22e+eMHe9QuqfwvInhEZsmQUqWarSDZEdor+E5d3lzJ7vCoDxi
zirOT2IF6nhjScTIaoIrA/bi8MpVYJeqRI/AFbX64/Ur0Ujvi9rUBim0FNqhZnBa5U1VkKj/Cnvs
UKCuTsgFZjnMdPsl5O03n49sQKsQFlsJNKeOG+xnRd7SuBGn3+//rDCNlCq0qoQSYidhQAUIfc95
GqB6ZGLtK0pP7rgBjW7gRowytzBN3fLrrclPDZ21cnoJl/5zoUp+6TLVG0I+XiXspI77Z7X5xqor
vfqIXehKKTl4AGNEIE6/xW4qZYMqM490jLBqydPajgjLmb3EOJvnEJPnzowDxgp1wUZw+jSNDNl8
IFWvER7SG+VQ5XjSUBY1qwbpXUp0mcixH9DfpksmoeWS5yekMU8DWbOgrDAKWzKLvbuBV6OY3h3O
ecrN/rw0uBYyPfOSOiFBZIXxf7USIKje7uY6wgy8hmu6Gkl84agyXR+RbkS72mSiP7koEEyfcG1H
3+RRjw6xe7UyC6zo8xrKjI9JQV2K/BEyGJQdEIvbMu/TQB3PxNpmbLA7HBG8XiBppPkCcqSvAK/Q
MAmKHCYAJ0bh/DIG3l51Y+rysKLC9YmNfOf8v5QB7Ovr7MlWDNQScwCq9eb8KQDC/xKEz9qgU40j
m/bmpP6VgnmJjLMaUzwiW1MmDIcPNwN21utZ7rbU4XGHmmvBrssLyvCEoX9qhWkMONMqNFUhNWjN
1JgJPm6B6atevtTaNuZ0c5DFIDaGLIRxV8qqM/53n9ASv+aDg9kbTQBlibztW+yVzXx6OsloONTf
KIuYkG4kXsHcYprxacZig9f2t1S5reb+q2BOYoiC00YpqqZuaGtqeRL2l3FngJuRzzsVMmmbNB8g
JzaVM6BuNuwpmO23vA8S8QdwXyppItGZ+ZecMLjlJ5jyW0P+MtzvjgXVZdOtrgRUmNi6UwqlVYqJ
HDKCr3hb1CsjdZGJgMF+lrqaHehymfGreUdoKx7Nk/8G8hnYgsQ25vwfPjAnuudueyuAIVWk/Cu2
ytZju9jEEP8IIp3Y/QF9ZxUUC64qbS1CrjXSYMe+xhVeeM2a2DpGxrE0cbHAj0feGiMYiCepFZP0
bOLEfGZkiNL9qFAlkxIWiOY8zZLuZObh0D44GRQa8yqOPBxCOxUz0V+wRTcEdzUW3vlsuAtjrtjc
EB0DtQizrIUspPtvtaQI7NwO4Dq5GxP32QEUBbV9Qan2MIoUAG6f+RgB3dkuEqw1P9jdh+mkA4CT
uwpzOeQ1WXI+pgZVIMDy3zIx62fFmyl+v0pn+yR/0aC06XijQXDYwnoL+7pc51dNiXNIsfl3A28u
UUKhzqvU+sLCjCGWUUjoC8WiWjvaFn2YEEvwCf3LbbsvPz1P6wcsQEH7FGog5Bp4PHrl6ZeI7zca
8dlRBu7wyE01SMLATOXD9JfH+8lMYd2kq5bewgtLaYzzXkELtcXkdpeFNl0vKKO4yUewEfidyUhb
lUzIGXjxtPQCs1fuc/zXjVzpcv2kMZvwe26RNWLoyxKc0Ul3PDW/lh7asx2HDFCGwqbvBDV9Lmz6
KdGJyGWmPDQAAEWRDWYTWgwoT6QtlAuIaP5xMthuDrnvK7swTb58LWzBkkhT16lGh7Np9TxKTEpS
IkcHsaDvXmljWi0TrLK7XmTGqADNlhfs4adJQ2irQpVGM4IlwmsOUJXO2cMxWzV5t4aJQXfi0rBP
fYaansWZ0GqUyG5KtcIHyzhTEvCpfcerSo8VSoEn/WBKMR/Mf55KRcCvvHHH5HDVimtsE9mzrQx2
ijP82uLhkZowE+z0o9bipvwbVDq/F+usIb9v4wVGYB5UM6tjoAs9vwThHuPDdLrnBrT8EZadXt1e
YiFKqI9A22P9EPvuZE9b02NXZkglw+ty9VLZlb7HZjIQhb2nPyou8NoUngggYD7cbIAC3AUuYBy/
0HylEnxJk6ENU52H3m+eB/c6M9efPXvgwabX3nsikkyxIferUebRAH0vk4o3mSLq9kJDQvedRAEU
SPNgUR3A6Gcqzn346/R3/3JXef9CMamn6Q8Nap8iTJI6BkC3GZ0+g/FjgbihEzqyXXKXkxn46KG9
f0TMtgC6v4Q+PxiKQtmtJQxmBThdmYobT/5TSB63mOSyfbxISdGR2eApuqu+34iTz7Dl1qioV1J2
InVQ5X/gvpy8EeT2C0jEhLkagGbXSrriGDKJnV2Y9KV6gxPop84X+UlHk9Da4fNNArlwNGFE/AZF
29cAnqNN83gDSH0BRZbzI9M7ivmhdeFvQ/xoQFHuQvf7IAmINsn3W6qpeyZ6HMAtlL6bx/NqFTh4
KhDp9e0yAPvQG5y70jZeP2zHL4v3kgSqFt/A4DT2Ni87QtqZeEkcrGLTtzjTBysBJs+BaOD56SXs
xIVSpokBtE0NAggLfggu8/cPWGyMnnxmrhSaeOys2Dkp8/d44qWABeixEBeI0nn/dg4t4lJoFzJf
qCfF96vJg/lCwFcA4PcrgES2SMpkIHWBZMnkE8UtiPu3voTmGSzbvnFPNGebegm4o608w2JidXdX
YexAKdwGmYYOBK85R8UQ+kDa+mrx8Ij3n15U2uYU0nnpx+aptn0OodeuvFm/aEKvQa83cqi5MyPK
SNvgr9ShYXp5eK0kT6E739/EMNWxnrBuuVc8A4DOMqDYA23VGcs26oXBmQYJpmk9lNgvrau//5q1
cjJOs+McuAbm/6gw7NQd09UOQQnli9uvd11NgPIFwrF7h6JDnuI3npRVqKvr/ZvrO7OV5yJwhhpc
fRJN6+J8e66LeBFNZkBDx4fZ2yOb7JBj1rQeAEgtse85G++L4IroKJEYp5EOPWuhehDceYMQu7kw
j57+jwPrIi4UHhZpx9xl8j7baZ7Zcff9dMffxg2KijijhFZqxF6O8yIoHVRJTA8ff1tHAkgZYRXl
Q1efxwnSWPZ8Jk6elbJVe1C78iFcfjMxmQLVlQRotJbEgFA99b3ynOtLXpKhpkzF9TiHhQkpabEJ
kpKmxNzoEiyDbuQZ8yYmPaf8UNRiMwlmRJ7psdXJxI2Qb4xmSHHw073BUWA8uvWs1m1IuwCenUYN
ZuF5LOAZ8h22Y1oafTcLYnUH1LPmqNkLX/loxqyVWDdhkNfHVP4CN4J5ibCSGEV4IoFS0ewRCQyN
88S9RAuhcpZp/u+zN2g7bOhMP+UtMWwHWAcFBz8oGNxJS5omt35bgEI/r0eN/sCVWjl3VVG5N9+1
WIcPLCPjtcPFJ6Zk2P56TeB5oYHYcJQgvvIOu0y4mXcb9LNgroOmXsGzOlaecDr1wISCuXeesBSR
aiQhU2CUt+rqppH6nnJUJWEyGkqAy9DWnzZnbVd1pM/SczokScqgS+y1lKvn2XEpH3KIswAVwySN
+agfBZQ5oBhkQ2ZO4L2qeYR1Et7tHYS3o1/IEw5RcGJn3HMQmjnX+R3DyxtMF1Na+Xhc9VRdomDn
Y47nAliItTbs0isTsPqyIjR60w7r7N7FyqaDoythAKMpfykXP8ApPYwTM4snrgFGdbq0JceZK02s
n0oaEzl0ZZAgUOSSSOH2YRuhLXsHC4XBufLAEau05PvSepdzJzntx82h7PJkS8Tor8FUrEVgTFA1
4zN+sQnnfdzRMVweRejWeIXxO8XFt64VJHsC4EtjV/Fa8bmMFEeqfXbqSOje05Wtx041FAdFCupD
XIiMScp7+AgD2g71k8tDIHGaJpISw63H/VPGl98c7U+z3H10qD6dYL6t9YjJPBpmn539h35ej3Cj
hyH8L2f3TiahEDNo4+Dq0srq2OvHudo8l2t6Ikqu4dvSTowcUPiKIxpogG+WnztFzV/cqFXE7RKX
W8gN9c+KzyvyHB1csA7kano+dfDTUeiB/dYf0doqWr4ykJzQSR8u1qiJ0BsuCcDTtrp8rWrE1bIo
7aoT86P5Wss2MwVaX2pcl6585FUoVQ0i/hV6nVGB9/oazZvrVipKfkoqWFYc/3zCthWRP5+KwZ7G
IT6XHUonQCozvwt0DqCedf0ocoTZrz4B9vhnpqsQrD31K0lL9RrHcS9R2Dpq/G+Q2LYYRBGz1Yqe
UZCGTPjem2YjqPCpOchP6r9jAhPz7iNQ4OTOMHXkghPbHSH/x1YA2gNREG7DHQCVA81D/PlJ6I9h
pNR94AzmiwFuaDgGIRaNMViQlZemYlguKptIDDDXp3hDw/Ku53iHzwKA5f+OPjIsnTAQMXfgPLaY
hP/QrX/Iwh/VnEUXuoWnW9MDTaKPANIaZdbV5sqbaAQyHKYPapCFWJ4NS73SpZZ5XQtwJQ5GC9Q3
HJ4xvoiqY8mXi1ebdDw4fYL5NRQpOyN4LZK7066FIjuXfPphxV9MpxqaBgMsfWukIc5nsoOfmSu/
aWx5UAbruUHkOymkvjCpGDjSUFb64ue2RIlb73G4rm3wlkzKSp0CxexBd3qcgzGff6Mk/i8el1Sj
/Jk6k1mu2ywfB412gYpSbYNmqssfrVaBwbl8p0agxEiobK4EJ4Ponqpb4LFL479zNePi+WIn1Bc6
CO7Cc203cahtpeymjeLIIJar31SkrtYyd0P2ROk5x//kV2KZ0kwpyoYM4hufnOCokidgjwqrlCdZ
dMo+xs67wnMHqOXRhHlGxJJeei+8kTXTqONHof+f/463yEPnyF3WVZgGpwLHTkh0Zd2tpsXdbuiS
08S2s5oM6L2rsKHH2ZiUD2vgs1PWnq38DWkOF3BOsRTbvuQE7+46IDDuaRZwnYvrXpqBETMVfyxd
CyuL2otuHy6XovKEHhVf/1ox1pZkhMSoBU/xdOS29r6Wda0SvqHQ+yxOfW2UJ1frEzFllnODqpPk
5HdrFB+GWbA35QRBUGoVB2h/HldZONJXxkuAaucmxRHz48o+5fu3RskiAG8kTQD8Km5f3RKSNr2a
TiGJYO05fgxzEtwe+IEExetBBS5Gx6SrjGubCVIuhuE5e95ns5a9FB9ragmJFfhR+HFJBO+wBf1E
tSRWrHtBPagEhLD1OnmXWh1LaxKpx/gxa1gzWGfFAkwBfDQqaUWeWNwzfW7s2pl6sPFyLwVun3bW
CFTkd7EUNhLs+8xfzT1rLKLUuyI8r4Xbj7sAHD0uVPPG7kbaoCwUEEGYb6LZ8kKdVMHqclsb1OQQ
pUAoVlI+wA32xbaZtqDG9ZSjK6+/efmgoXmsS5pywjQ+H2QhWXTqshSg08+DjCeys16Kwv5JaU1+
aR0otfawHicrWfnDM7wVNT5FoczZgEeUviaLTDfsdPUEpQTQQiXyQkgcKftRDXRnsDYwIlNJdYcP
0ICGi8GbSoo4FLm44NiHSILn3L3X+IGjZOO6whuG3ji8oEPE840bxXBcSteE4Mfv+yJ+9yG3g2i1
RC1gDtqZb3rX8P1uhCLQhHTzSu02bRifj+1TxJ8iFh6S76d+WIcEiUplG+52RNxcNRbQLVOePC+g
8feukSTQwbvY0qxDif/+rwuJyPTI64yBGaOz577KwHX0Rm/gVGrcL5M4uxDlF/PowEE4xOM+Mong
k8r4RHZWQUv4Eh8cLjyUwnrHGip0LUn4vvso1LFTRhfdOZIigH2W6XkKjzbmsCpm1frHQwVt52Sr
Rz3t4yxxmmbJQPov+LUk2WgHhcHMN19dcHH2a+vUetWzCjIbyt6VmxqOkiueuVhhqsFKwSWw++vt
YvLOwXL9FGnHu6SepTgwzDoNtCvSdNUK7JI8ouuOxn4jY9dbAXTRQNFDLzLivJarUI7D+Ie1wRy5
aRc5G9xYjMaYVU+K2tQU0qAgcT4/Zb3RDHDz+79BvkQ5WcsR6sJeaBG1flrDD2n12Qy4PZ6UZG7o
Bm18u2yuiAs6GiWbKnGp3xrltqstCfYuSX40PGH7lpzBGoPt0OwlwSMuatSR/XOYVNcKWeCtLDtO
DU2+2eBpm/LQB9XkMLHfMuogTWag7lw3MJdIPPj97VUoB9vxhSJlieE5gIWzZmdIKoA5DLmOD+zB
IUkY4g1fIF4k69fRv6Em/K8hSTwK0AAXd08/O1qCgBnsZJgad4KprKB0hC6gy/uE9GZqfZyVFDwM
30+tvRix2V0Y3XSBS3imAtaq0BZ6nrBU2U/EQq/pT3FTqjY8iKC5Wks1TWJq+KJYKuQes8x2gP8T
lGSoaMSBk+fYJPQVGYCdjbGE50MWHGDToFA20YeFGK3tJnh/XNnrQ+cI4w/aOA/yc1wJsIla0qh3
K7Hw3PdIW5GLZ/1UbtMNsEJGux8nbg8Ae9FqwxGavva+k6x/h4Ifyz+lern1vLhaWFB9bW746Ea/
UEMFwxbNJ2Nm/0FoN3AVP/vRZqrPrn3zXF6EK9rMs9JV7NLUWFuInYn/odZOKLW7iBicIp091lKV
OJbdXl46GLigCyhut8a4OyCRD0YfRjXFDMMgmajRwf35yQg1HrMzUkmjVG7OucRSX86HKBmnvoER
zxruvvTE3VammjXJpurtalTvXhBlpdvJXFOa5ca/KXzzTz7RnPrXkUTRKO7O6NnO/WqAP7O/iyTr
utK0ClmMLU4xB66bN/sD3HCE5cl9b8z+GNy6N+7zDS7D7wPS6JzyRIjHTFSTlRFBQA0dyPCqy7W1
tlU9KkQF81Uj8+zHI8ZtWEWWNuTep5+DcFHxyoWwOyVUqd9/VG55Y9YuhxRWvlSMs/kDxGyYh6n7
/b0j097mctpSMUZIrl22ba+4zqhQDaWEDkVgJRUXDTps2zyflfU+s+NarU/RDqqIZeLKDr+FcdY5
Gh/fG2LRtsAxrFVAwj4vdl4Elrf+b7UJrqQDI5PQXoFtBylaomX4fWJJgztYcV/NFSVTROhSc4tE
enU8P8s1etYTosEMXaW3fziTtiYLG8yV107Eq1rPjf6Ml5CxzNOzihNeed9BeUdmH01MMargqNVs
Ik86QuYVheURjlPs3/lsxhzKPwR+KfAMmkDrvIASZPZj35BA6LT8GPcZGtLtvPRG8KV8aladOpW2
fj+vIpzQauNWb/ElG7DbTPNI/BSZG5fy/cwcfrUBmHvvu4Cpdwk8o/Ct44fBVeDRdw7mx8QOuA9b
kWXPiO1GRxZnEUQm22UwAGiBv/8XV0VJHas+F/SZc2PZqMd62zAWE+klKehVlUZiPEdOIZAGE7Bu
n3PNxinMl4K5HjgHci620reCvOREleeWGiOs5BMVLN8XhZLm9uNoRbya4aR38BZZsombBB7XGhf4
/riqCF8Ivzb9rQKa+ouuZuX4dHDG1WLgjKsKa8pJY8IskCjtiGCh7ld/j6Gf8vDz0840c1tu+0i6
5mn1EMmN7PI3VzwxwkhRLsi+Ij2WEfh8Mc2AvCvHiApkMAkVitExLiChfvmSVXAmWyMQSo31VJU+
nrmy/Wu7MJHDA4UFaxYfnqayompM2MFcS0tk14lYG3mP0HgqrP8KD8yzd7rkn84C5j0CytgjAXpb
/mQ58jnPMDyA/vMvCYmJs6+4RwoL4TJiHfdyiXj+K8rfqomMThRLH7KY5T34I2sJwsph72RJBlBu
zx/9sN1q5KoPBo0BRsvFTAhOUKHsMQ8Viaq6+mp5E1v+luyE1F0HkZO1coy4vTRI1sEI2JA1+x8R
SvtQToqHfdo5PbfT9oDdWVmtioGnDg+2MIuLAN40RccCFVuDrP6GQFk4/QKNDTqT/VoekJe7OZb8
sDE5VB+tyk3ZgXgN1k80irZyG7rhRpeK9QHa8iYUX/mW/zsA46xbxfG1xfONYWgUK6v/6ZH57n3B
8dFH3tVJ51eDBNhbz54PGloX5Wvhsv/E57RdgoEzxga5o2CIdwcWj1ykZkjfkobGQTUeBWEPjwtS
nRE9unKzv2n76dyFhVRrvJpn5H8+ePPBZGrTazTHYM3ODZpUs1TEixyaT8u1L4JAPLvRLkFuhEJ8
Th+jaNiazDdgn7R7UMxOTB2MQw4x95j2YwbFS8wIfvFILfXtzXPVM+m6BZOXRObRCB8LU8LrsOSg
h3cQG0bt0E8t9MqkYSh6nYXrtdqB80EwClxgXilcqGrtzFDP/rRSHpDff4DHVWeTF/MQC+Z57LDw
IN4wRc1H3Qqd2rzb6qZ71oeI8L/QqU595NmnuJbj6WD2qAkrgWqY82nKGbPSozBTVywqlu6STSMF
eSIhajfxma/F0n5VYfbrne6RgoRF5dhcw0LMlY1Kr195PlIfaQj57xX+1Len6nocQTsA3C9WcRBK
yBqz4JkeYZ11aMymlLnXIh61rluNR9JM21tLTmfUXWez2iUB0uWNukYmyJMTbIQN3fUI/9cZSSm9
B0su1+cyws88EN+nPmbcKSYTLMqjE2S29jZPGNWe59bGT6f6uX7BqBtz46fRa74BwdXYGuWkVJP7
aQBghu1j0aSP51GOxV9yZy4TU4RbwnLhc+ZAWnEBZLEWi8IsCwjhG+1n6KcJqX9S7HO1pRqYjpxc
PjXqdfW9A8qzxwhizDs6TvC1kqz/gwGbTtPmEi9Q/4aYip62G/v/S0E4kdjICaxXJ33IS9mO8vli
Pl4SonxCNPzL8CyDdbQbCEO4dSFMHXph/6eAEq4FNcd6TbAfpnHscbasq7OMtjrQD91BooLHdLKR
FqrR8ikpLQml5L5zJi/DAchRHybUkGmvEPSx54QXkuERImJOqNmHS9UAcQ61HJSbraPzFJQyNBRF
72CA7w2AHXayq7K31/MuDuBwo5z+JUtlKhvF0ae+NW3HjRSYdal1OHKzySCgDesaZhMyl09xLT3d
AOHLLiahhLZytcvK+OeJCAGD8KpPvL0cgwFgn4FMCEkBw2or6eNWK69aCSOPd+DgqqxYK0h2EtEA
nvqY2PcId0mnbGdwY1/JaaF97nFOvKTr9IBOsfCFfSdQ3iRozM4eobDhwIQzjsF0HzkjAP7N8cTo
uH6475GlbaY3KlpX5VJuMvkczH6JhCZoW9WV9sPNkWVPHw7TlkyQDXlld8CrvQfbcrzg0iU0jhrI
jr6v3ONnC9iqd+YxzIprLbojxSkHHoDi7rFEaTN7SWhbbpAdD1uBhwty5aG1yuRk7NgPQDPFfZpA
yF6y+6gY6Krhe8kA3knJoYO+MPr+H7bAYL/A2YlxSxtsQUXjC0NVNyzcSiLhki8uymFAq84v0UI+
3YAVquFgy7Y0+WF2wKSzK937o/O0NnwFF0uVYUGzzPZJrgQI9sNMAPEtugwOfpi/EWJbbXd13L1w
2weF38t71ADXu9WOesoFIL3M+F3NrZhVud5ekLFwy5QJgkApWAil1q7ZDxKcCP+c1kP+WWfRndYh
5dCRdvUGaPptai7InZK17oGS2KFj5994Xw211ITebIqtSdE5xNkE+/MeWMSQdLzgHC7kWIjCZz/S
7qLPW6AdiKq8JMC4Qp6v6SwfaeT29ExdamPVUt7uVqfFrTIX8SotQnUgq7bbWZRPR9CXITrBRks/
0O4NMJ6EmmkpkqJwjiEFDZwSDDgOuF5coL0OUPtyr5XpdBfaiTTOs8JnRQ4WdXYoteu+z/mkZOn2
N/PjW5kOGa6Iq05VD6IPadIyjLdNKk3qlVpL9JZd3BNBRrT3lYkHsFfxpszeSqfIz4L6ZwsAxO8Q
QyEhfZ0fPow4XxNTf7feQKzrrxeA1Zde9b84+5hCKzGUCRS4zjaxCVhBMiDGzSC2R+a6mp5aRQu3
Ujr/TwEoXpnh7j1L3QypKv3htfK/T89JMsX8HnPFk5dr9sPIN7PDkxflBLP2vBbBmeMYDtDbHMGT
3nKQ+d/2x8DyNH7fwInxFOtU0uayi/v/BQ9Hsh6nPwzxEIjQ4Sl/7t87c59RQFMq6FgdlqyDYoWA
fxczMUE+rPDFLbFNmyr/zdWZNJqXcgiigS6dkMgCs+AKxLxh9bhHetQX1OUdSVfFIGNBu7kCkdAh
E43CZnfh4P4Y3hOaOv8tIbvZMM/sX3qJDDMB7wxOKuteenLlM2A64ugrYUuD+7+HApI10DrS3MfS
MPc01rjGt/9oCcWPL+RRSI+Go2y4woHayY2A7E6xxJgA/Qo0I98I+kTNo7A9GywRv8HQ67K3MZhi
bm9HbEvlBs21E7pRaBuI+mB4VZ0Lmt0mhqPzxHpvZqwm9gNLRXa0WAYSKOLldStXckCEd5FLh/yf
LcSGMoJZIs/ZXjjQBvDKKdSvXfXrSWfWM4LNdBaiRYZU446gms7xYgSR9bJ6p9HrOf1n2+vW2ili
GVHd5c6oRJRrqDCuEVoo3qyPII+haM6SN7irEvhzdgWz2JiYInmSReyAeTOZ23yovhYVTXBQGLUS
ktSEjkD5JMVKvM4+8NwwIDT+eyGrWFs6KNYQ0Q7Uh4TC1k0RCOcuSTDpA415ZxqW5hp+SOfhvnxj
beuahhdBdDg1a+aCOUnBYYZWMa9lsnpAkrYcLQNxRJa/mudyP+iTjJK4cBUpaiN02ObwDfqTc/I4
hav1YrjhjUQLfbeLoUuYZxXndLzNi+1D2rLdFuMnGyBlDhN5JCihqSzGsoLhemdQK+fCCi3B1qdz
AY6or/iCYz36X/P7upAWzY7Zsdbuw/kuvqgxolktFs3JHOB1ULR7105rVrUrGZjF5Ow+LsHkf9xS
kRbLZtIYcXVpyMGnJMpc/lPgvHocGzccb2kve9XmGsnchn1dE7wGAGQmxQGDHasMMH6SxE1f95JA
tJFEDvJJ5w/kF1tmkRwE0Bm5JQGGQDvxucx+guS6vQgp368P1k8ysbK4Cqyxv7fGdlu84rotlzcI
DGoNUb7liBWxUD1fABJ30VhBwj+jlx9SBh23ohwhv+A1O/RbTLm5SP2NzgWJWx0lFB7DAq8v9A0l
P+od7e1wP55QWPeHVTsLInUAdIdxlz4sbcSvWcBZcoTm777AZgm9DE861EulOHKC+0N/jjnCGFg8
Y+U1ndyvGNcTp2tgTZJAMZ6OXplOLqeDZkClPADOiMie2vy7D22EwXlsPO4lVGWnZfParB/eCUes
OSD3Hz4p7eazZJ+yczzsGTTB0D7YS7licDZ+IMmDVgnNA2d84sLjREvNyjEPlHpJj+o6mMBvUkZC
Z4lou6dKBdt/HA5W2iKcAdj74OOrM5MVPJlX0hRNqqMFN6UvXUc08E4N4V+VXbYTaVJO1f2NFuL7
CKbQuNjozhCUKHo39HOUJ9otaaWsaA2koJEQuTPzkVijU4Wd3mbp/uEpo8j+bFiLtSqExPAv7rNW
n4iU18diSksLsPC2Hy1h9XVvkIj0UmkXym0fJzdlCSzarCTOuYKN/PIaCUXaabua6v18ZIR7Tyza
9kWJPg+ZeEXTIeT1w1+GxM+LsGrfPLEyK3d1201/1KNvsP2ID1olEp2F90gbaeaDyeQOxBUrYmpO
6O7/Ng/eTpaM1HR5HKh8lnYxj3Zoanx9cl+O6tC+6s1O4YgvUkfbVcqN3XWSXioD915WRphLk+zL
qweKrZn5fQOSdM40TB0t4XhnksYuagp9po0QZ8LJCdwyqgtchhTRcJx8hYK2g904/FznVH5RoGwK
RmJwz24FXWJJIMzHpbRnMftkJoaJasjBVfdO7/bNd0Lh1LC+B+vJIeSOmsXdqbymnGpwhIIt+CjF
MRGnSiiGAHOGogdggCFKr3Y0QT5i343vw1qkuREKBAYhZjjYGmqDxxZGYwOwSQMI/NVuH1li8CdY
EhrZ7jiD/BC1HHMp6EBDk1BPNE+JC+UHLnoWjc9YSNGObepg+YinYW7EzdJKjD4KSh0eopXJ2BOy
+dMytnsDyAJBGS04FbQj3cxQXfupr0jjcXyRtL8dAnaTrLJVBeUNsIlsdDe84ZKzVEOrZv51Ql9h
LBkEjD0vNeoW05MDZ5JFBKXX9d82IeKlyxJ8M83ei+2EW5uGKGLOsmyK9BW7T7lWWUappDQjrYEb
fm75OpWXdqDdbbIL6vgb1VAHtjo2lhTlo6okYqT8GQ4VradizdLN8YBB0+m0N6JRb93DeWBPEFKI
ZnQ+O7pivL022q4igK6S7a1nG/qijUTQxw8zzlnPW6cVOQy6oSKRP6baKn8TXmOc/Bikabbg41IJ
nqQb7V+wHk6DJjHB5S/bGnb9bcazePp6jRRWzzaFnT8ajKgyL8WA+QyiL1EFqicDRR62lsENW+Je
CPFQJWmlGOUdHGj03DCAmni9lU0p9cK4kr0MqUCBol5PmQ3jvKWOnjS3/T3ElCaryWp2pEaY1goT
y/CfJ/NcuiVwbr0YZyc6IM6gsyIojLbZuhwbZu6g/iyHCAO9488rH4u5wbs9e7ga5hJEbDxpOnh/
0VatfztsZMm1eA9qX6KUGf2G8RVUjgkqCEjnVYs7Q2XRCSNFkJZ1LHVC66aAbpE2DCd7sA3kW3h8
K+sr9g1bw9IbWkzOxvimbaIdxDMnheQCHgWvV17SrRemnix4ythq2UAYwbThcx7PsvJaWRUZOuTN
9Hcq2CVAMIcErHQ/Ief7MhwW1IsNSJVqlaFeOfRzF1/AU+Io4k0SKCSs5WNKiF49x/BIVFkFQRoW
dnGGgLU9KBCYnKrWV49NNv0WneLY2k88K3OgV8E8qSkj+4T31UMy6YK69Hg7LAtB24wY2A6Lkv2n
1/xGZZVyHY4Lh/eI6G7osKjawf/wB/ZXTceUuCsGqArF/fuiQD1gQ3ayBlm2OLq7vpsxh2bH777k
/h9CPB4AzO1wYqMclOoYnRx4QDurHTWHR2U3QOxIPPNAp6QMCxXBFrrPEyyDXCOHn95fER6/O2Gv
3CIDHITHv421USm0Tf0i4Uxhi8i4sv93rBFMjrhnacBYOwT9uQAESBcA2nTxhO3l6KTZ+ikLv5My
fEZDUycGru7pdCYCrAg4xrIwLcRpFtB8AkIndiODIodsj7gGSMs/HDjbFKETxBvv/uhGyOAqwqN5
wP9a87YCJqDr3IrUYcav04DJv/B2IF77mkpR02Vaa3prDpdWlTkSqTW3GbFSW6CwyzVQ88Wa9LH0
h1CPj9lCSl1wGWgGWXY8f6vftXZMVG/yzi0FidpweW0SnE4EOcKacTfcJ/AdyvM8UHCpZW7SL8QR
CbKHF5lFTXaDbUoXwGO6T0OUuUf3h8F8OeCY5TtB9b4S6IetVfH1p6rvcKjHOtLzScENgerf8Nfw
1pJ174ptZB0KVXQYKo3IF7j2YTn5M+pOBLGN4WHx2/8DYHg3C5RhQntlIPLkKt69bpK1lBwcVOkE
g2jgdPQS9nyuP9F8UKatPmSr/jttaVwD/Pw7iUi4mKzbZQP+9+c15YPW2EtV5VDRcM+wXm7pROfZ
63rpY10Es17C/DplqIwSHxRS8AcKeuofBtxnchj31wqrPtucT94zyHeuk6qG3IVfFjrq98HyTEf3
5Iyt+eX6cHad4qVff3p3ZdPcvdWv/+L9dhdmgSih0hYstzw0VYO+miHT1/wElG6jeydpogF8KzxU
dXF59kmGlB2Pa3i4NiAfaqlrLzvY/pG6Etagmb7TgO7xphKehTl130k7P62ZY6XfblZNNZlTyk8E
mS3fH36+1LwQG1G2aRXZsCMEzPfZUUFGtULt0JkXf2IIBZ2JqtPf2aK2DbnznPOunUW9yMIEBufG
mXabgkp29BKkD+6GUUkWIIZkGKFNHmQ2hvzuq3n4ykNwVnWHxIQnLZJVxqJcQopfgRbY64ir1Ogr
QFPXj1xHv6VDH+l8YrJ41RL+StJuVc4ZMHivsSIMHpFu6iE7mcc16kVrGUkWZD9nVs+lIII0lfSL
GGhGYBkUQJC22bO7U8yZzR7Zg4wCoWDEnhbZLqBxvfOlzk5I+b2aaU7iQ2ZoABul5wnR1cMDw+xB
yCUVFHfXY2K1NEiErvTDURn2eKu6cC8cvJJHtHCtWyvWKkVlyKZQgn3EWRRhexzrd4k1ei3Y0/i0
YFbCxseBfecnRzZx/a71q0HkqhvxMWDIamL5g+/EIUvdEZ/ax3dmOk42jLqr7RY+mQaSNYBRRNDd
HV0ax/4CaJ/uimK057roes+xfmEs/gWmWpuoXYy7zZjTZ9LHaePhrlAOL1V6VJCkhR79Cmj+F7ZU
BpUcTCqTAhLyPL4JSr+0BaRzOhY4zOMzOUxssRk3/0+Xxz9STjwgYjrfpwtu7/qWY0cSnoFP88Ku
MIeZtw1nEXs/LLSYSuXFk3iZ/wtYgp8wpYe3z9PQqXPO5HzDQTWdEmgCDZuUBLCm1r+tkWtjRQav
kqIx+pr1Mxr6OdbsP4C87hzwab/OmtRY2niSSPM0m9hoCtFOnw4+p8VN7GZN7lwqYQn3HlUQBla+
m43fATzSzHXl8ph/MuuM/6DJcj0uOLKlLISt2fbQSV7b8zioHovEzOLMzILM5Eln1/fu3Xqrrhit
i+h0+nrcx6QNN0inKqotKkHYYhXLey0hv3cRCJWPk9h62M/Ru6jRRWjjse0B876wnbh5xgGdcesR
KQiSodfRdmFHmjmuDB5L3GUwh5AzlnG+fRaVfI8eUVcMStcCY+m4429AS7XbRZZ5J4x8eGpMq/aG
c4seYkWDZuaNwgv3uEhFzfV7TtJy8OJ5MynF3gpkK7LnX85jvb9B9vGTvzIDqA779ViFTYnWbXcQ
MVxknCvtNaVOYpWezrnOiiN7PBnRm9l4rilvdQVKxGd+22IDVplE6cEzDXZdI4fUn9Wug/4R5Agc
dmGgTqPa5ZCVjxkLA5hTXaSq3HU2fRXcn0fZ3pTwyadJ5Wg8hFw9tpYsLsKwVlfo6f9TadVBXKJE
z6OlcsBfrP0o8frz6TjNk84ogdArsk0jQP3UxXQzh4ltwGGx4upS0m27MMOQUABb716qIknKfYIy
/8cmEGzjqB6PmNN7qPHm58fkEDNKc4AqO8TWGWg1d8/a8Xqjl11cytasGzpRcfGLugErWFiuG2Ni
ot9DcREZB7953WQDWWTJFD52AHytFbemY7/o2Sqj5osXrEysiUDp5EEfwVIim7bbNkFK4MoVz6nh
joBS1WXPjcKKpTCRCMZvtLM9o5jXGZVAi0OPZNlL0r7HpV3jWXkf4I0OPd/NS7JMplQh5lYu+LHt
QkZoLIDnUrh/ZVhJgazyDaUqjvoRf9lLmOJa9p+lkhp+GTG3FuyiXJA+XuXi/BPQ44UjjBAB5ayK
P7sn0fbhvUZZZyIxaQaF5kjFwgpYcmrdokFXs69eeSeFwYDEuz/ZEaGqUdeL5QtisKCEzGro2gx/
Rt4mRm3cCa8YiyJAkwdqLPSiTwerv+53bh0l3Dzx85QRcJq2fsX3FeXJ8Xetib94R65ATYEX0SZr
C8V+Qc58IK+jdy4971AXrIRnM0hhwTrA+/VXINpcuLB0MmII4yBlvRQH+peVrQUMCyUov/X/reL0
Ynd//W3m7EKPrwQu9vVZMgYJpIat2FAgBtDzQbZ5VOTj09qpsNxAeMw66osiQpx8Ryx48U+xIx7C
V4ZdtIs+VRK9AaEQDNRgW2F2wEtRrjb3a54WwMp1lnUuV5jYVfVL4QTljNUsA0Pxjj6x+OMAl16c
ctb7MFDs2BEpczeSUKAr8C84M4XwrGcRRbC4ZvDVR3nz2zVplPKJ/2o+c2LFfMrkiZdHgmqdxjW+
WBTtpdvg1+QvRcmljw2+bZyITvivFzsd2RAlZKqIXqi5zP4njvTRhlZBtVQRhpYpIXS9mFWPmv95
M6M+HFV6Qd4y7EP6LsGI4kKYFJe/rKrPqXE2uzRWY7yCti19xizV6w7JDL04hVd9zIu24P/gIWd/
DzkCnatoZioWh5E2Nd6M6QhghNtJAt/e1Knz8K0p+07VNUcz4jn43hFZ3IA0IvO9/Ksy9pDxhMMT
PtuCbQET3hNEfCEEFYhe4hmvypl31PlGHMPjCpSVzIgZaLU3cK8MYw/G8rzlTtkqiXNbcOsnKWZb
pP6/qIRikPc4Bf14STniyjLB8GVxqROf3rr6S66Joo5n8JdPTa5BB8gfUEefV3nTYBIItEKHtntA
JXNGTHzSxyfszINpCuoJrWqMuxx1KGDhgugh9K7gVuSrRYWJthDzAqhgporeZMPn5+DGkY1RnRvv
Gu8x8/iY4ZaRJILOrf1zFhtH0SunEY0gTYSGwrTS+JU2D21tsutm+81Cys9L+gC8u5Q+Q3gmlLPF
MWctQdpB4mrfaANfuFgP6LGGKeGJMBg372d5MY4AKhvJMmVn99CSxvIGm7KqHT+QT9Vc+Ib9cw0O
WL5gKeySmLstC6tBDuo5r6W45IKNDKRd2MdqIVlpeS/uOPa2pfL2D0HGbmGvfSbypEjaF9M4bSKT
6DUT1IJLsgJrOnVT0xEv25pSo9IQATjDM5jZMBBSkcMce3NWIhuo5KAXNI9d8ZSTWLaPFIAb6MC3
YHdDKo6OzYGEWsQ5Z9XHztdRSjmln81+Ohdgb4a0mnN7H/vcrBXFnYKy04zNfgcLQEKUUOixcuY4
g8BfsnVAQ0SbgOIWhObQCB24ii1Voodq5/3GnZbMaVKJrpgOMUmnL8uP21xvzibWx6CkFKITesWn
ZPHPzpgiShiIw2SXhauVW6lGg1LsEqvxJsUQ2wDVRBsyOXJBF6fvKa4o11i+bRbqZvMzEoNcclvE
hP6/f9jht0a90RYkLGG1o6cqmrIHXySuWOnOzKo7XwF/aFCpt6nCHIfbqN90yZQDJzKtuuLO5981
dnA9+5/tMi2ggtQpL5eWlnzr9xyTKBw9o7Sc/dMpWSlOxpx1ES4CbD9Ts4gj6nywwlSmYFEoaweN
v0GoYCwkl0YWJSKbvnk+K7YhZB8sgs5uonuYM2nw+fx8TX1a52KuG1HKh0Wnnk4q1nyTJIZzxMLf
R82MP1zzQTM9/GKP23rcHzJsH/+ebr/7F5kh5dVpxiDKcdpAfPXCJBXtktyc55VdosTo7KFpYUli
uun+xBwMe4BeHFBhUZ7hVOXzjWDOeRk6o+f+dTQYKIO87v/RB/ypnCs6pmRPwQTA22ItwiQo4hgY
ieHpedvgpH+jqFgxknFbH8/+hCLH3RRM0tuou2pRcl04J8vNHj0577AhiO9ThXCIbTYbE01IPO8J
Kx/oVcotpV2XWYPUEGhzlJi2+LAHNILLDlbkTue18hOShvAZ+5v0VvBeS1PGDvhZq71KU2sDW+oZ
nL8RsbY/j6cwcPNCwIBnCtduUXBzf19Ng3rZZczkFXb/sVt3u3KueIzkGZtbYmrwSw/m1lBjWCT8
zWn7BvtQHCghUk/C4v3lCl132Nr4I8WCToDO0K22MSb0TeqLRojWTaMPvFltNqS3Ao1Aid9m07+q
gY+q1DakgQAnUezKKlON5uEF/kaW7pJUxRhAkFe6CzIbmPS2wVEHr3LNKkdaff/ndHafqp/TJi5v
rknw2D353d1PRYcdxT2iuC4VeYBSeUVEuXljUPZ7oB0BjA+9vmeT6jz8rmKKkhEpG0AeGh3txydK
H6Oe6RrSMllhmoZ4i4Ea2R2OZ3kmdG7pbpNgR6OJ2mym5uEwdvr4vxUTRG25UvbknwixZQ7DORjj
O05pagFv/TOFeUN3OGuhC5zj2fgG/thTpmVnRONEI+Zs4U1gi0zEzYfiwT1eDTnaYKLneXxLP8CF
mZXjKBNjoUTZaOtfNKV3NV9XKFKicDsGzlTqW4tffBlOm22qUBLj9evF19MRLH0Y6fPWPhmi0Fpo
4/9ra9T+lHMsKjWKShAIwQ2RWPg4+YW0ZDqfqa+V2pIq2KT2WAwUg2OP1aSisUPL4f362RgcLsQQ
IWE1aIQr/7qH1mS9iapVN17zwfLxhSlomnyl7iMDY17MdsJRo4+NcW6cdcI8lw32/NecqQL0ojys
bWTu45AoiztBRmXxyY0VZtjsTmxLa+mf1WVx04K0dKAOsymIrxrlFiHkfavtRj03j7OdOenVmgFp
6FMtekqHiWaNVyrZz9z5aAwWa+Wy5H/UDuiZ5S6lU8BY9a1ojtn23NcWE9D2zZEoiMTFTqG8r3vE
dTCEUVyq9g5IInQO8lUXjNv7gw9Coot2KUV2adS8U/OLJZFIAr20BkqchLQIZjg3YXgsUI5iTHUE
qP5XLEdP3vn8/HPGANWlVTNeoqjYHeCOwTEySPsRYLbTAdGc+ds3I/JDrR6zstmHz+ieRKgnfBRq
QoPlCxDRvfO8yh/k7mGLiQ/0jK/2FxxOKfp2B8cL/OwseqGNBwCqiwTYi3ZzGU10xCZc6WjwI0Lm
/9HH3zGw97jgEqtQHGpvWsOm0obkPzFoNlR8w0+iENgSy/mmJYQrCYM1rd+M6Hrio3f/9B8CjKb9
A9lrekRwQrp6hsijA6yJDRC1Ot0zxdvByaUxo1jFXW2mDQZGMms1aZHhpqXjCHJ0POVbXcf1uAv2
Zc2fABRExQtVBUXtssGSpZWD0YPEZqGEnbg4K2XayTL7bfPKZKzm1VP1Me9rYYq4GV/qvTBvV6Ow
gogQMqI5lPRXrSX3l7hXl6NGtKZnUzLHpKSIwwWIUZ0AuoCLvL0oZc/U6JHsxoT05VUvr9l5FW2d
0AmuNvLxu2IpVJViirVOwa012ySovA1v6Xjq67PE9TqEkQ3wcq04/Vg98QSGzc/4rlxQ5UyiOX7Q
ZomvawLHgaHLxJ7OuX51TSDV2BsRYpNQoNevrJfCGYXxsUkU/lFOhC0C3tqzn3h+xxby7rCg4jQS
x5HYSvtcYK9ZkVVmCaMkDX/3dXRA4SDbUNMqRpUn7OkNY+ccEVCqh7U/iVinnI++uFTwfDjBJ+wX
wcWDuLJ3fjfAkTsQDqQyXJvskenQ31cDzAxGP6XK/etKUWs0nc2wuyfx4oalpKIV4P7dgf1iAzTv
YLr6VJz+swyxqWKj2qqtLC6GSQfWnC16jWtH+OSsFa/to204NCzvCEZUSb4x0JMgeXxIaXAbLLw+
DOdEP0Cl6PHzjgJiKZUwg1dwunXm268UXeFun7tFUCqLz0TQoTtZy89LDSqGJmF/5f8TA/lg49Te
0zWUOX14K4u0sDYYdu/oNQjY/1MrvMi87xgM0vQ9775wVfGQqAqqkY+AqBfo6d6lxdK2TRaFA1pG
HC876Oipof72tVULtLquiAWkugtCNeAB2eXff9HXpEE8n0W7WyQ8XpUgfV7DOwoBRY/byApEDDJV
jEp4CCy7ShWuW/71yu3y+06/0KthEcx/oNbGWdSuoKfPFPjVQJJWd3rL6fgkfo7xVG+WesS1PzK/
xdOTIn+gIJgp5hh9EBu4/N3H7eK8AdqRpyOBL5Zo3rMq/3y6NmglaOPr9fe0oW9X7Qx3hmqJj8Lt
bmfUZDPt4DstKylpUXn5CpSoQkIvoA8A/tQ7jz0EHOgfi3R+/+2AW7sOJtEJMr4OMq08e5x1tHce
IOgky9VKjYJRbDIR2N+4xQ99k/iodMJ2xkcB6i25uZVj7sA/smBGyTcGnC/P9htyf0SID/a1+SrM
IceRBFr9JRLympzDunqGALBQdfC+Y9N9t6ZCPdrs/nXDUv9NftETnNyMlYHqyFfNtEv1GmXBpkkb
fXb3WQ8tDotKgP11+HAn+OGpRbk+WWiClVtK5ek83wmdQyzzF35vV8UJijRacp4paFZ7bI5YccJ/
QvKsJMp7KBgmuZoj7VkM+3Al+N3Ln5PhjxlirHrfGk+E9Z/bZnxVXQsH47yggupGdFdE3Jc7v3Tl
IP+vNmkMFSWtQuAP764sg+XqufuBGc/2sWhK5YcRuIq7XHNkGlAOuZNr/cjMykRIrmPtrmEWsY/7
2CxkqXCeRdggGPkQGS7OFTG3rc1XbiqPy/lUVF2O5s6lr8fHD3QD0+k3l3rFdOLaDnroJFLFiCoh
BNfxIfO0uhz/K4P6zaUBE6+PmLVvszK6E0RUoFjn6h7Tlzp9fpoY1BCp3ywtvP+LKAAAnNX7XVNO
8mur9SdktRd1JEyQgJ7CJ1RrCJftcYvr3jnhDmm7tMjhYcxqahAE2dqBD5Yx/EqzgNM9ieGvIhsz
RGxna3EKjSu2aGdtX8Y7aEi/WkHEPWcezyTm00OPsHa1DnQYG6DT38Zo3pUIMzK/wV1K0SQh3z7z
wMIP1CvinILldRfLOOlCInuhchD+g+wzMfFINz6SSZ8lCyJhgZDSM/4oN38AriUkte0oNLJ7qb94
fWHRn26fB8OazC9vTwe/BnyztDkLbo3Ikgtk8n+HXUnOl271LX3sK1SPpx0Nh09MhFq6Np4uV9Fx
hByBa+5PJnk6P8cwjkfik7sq2ZcgKrzV38KcGUBc0S/4v7mAm+5i38GaeCRJfEzPKgiqt2Btyf65
yHJQ2WxOEWSAXrUtucSZGTnQpxfsAq4GYrKH6+8SX+4osJtQPhRjLWRPwEUjgPHVHmP1w+2VOvhG
3qTwHe/5l2Gm31LVnfdef7lK6ka/CqcvSdCv99WvpkJm0p5ayLz/EEQ+x/bLPbShPKSIuN6lCJFX
PCAe91vjlCW902nIUgBt+fw/ou55KlkE1atqrJCENBHhUTvByYNIAQjBQU1NgP78NFLyFvH6rbz+
wx1D1bwvwmVI4UIRy0LspgO/HoTCf9TOoPjzcATrTGNjJuV+Fxz4xk3FRwM64OOi6K66mG17n/MW
zV5W2tRTwch2+WKInjhpuOimqAfCIw5WraEpK3UZnwPgnpNVvP++wQinN7YiohndZc8Abz4pScsi
xDPWZaHQ9CFOhixs3YHyrIvnHf1Jk0q+LB2p9ibt+ebTuP74mTmbkAFWwDC27NnD9zsXpTuXeRH0
nwsImR0hxa1kEUUEqcQUpIdXjMqaQcZ//6tB5tiElNdIcOcul9F1Y51I+pAGr1VjBxCDEwx8NcOC
6ojef8Ml7mwmL6DEUPoMqhuoQXEh5ecv/w+4x69K2ZDBkVOo1vA9juHKrdeM1JWFxBe4QIUz0bFY
LS5rKDtKE1mJ8fJpNffp/UsZlUH973eRCEh3Vjs+6kc+PbzP5xCVITyCJobH9Bq84RULr5XqXuuX
En4TlFqxJ5d5vx+agdHUScrwkNxKfEJfGBm1jyhF0fBqWJd6mNjcGTVhbb7JH1jPW5noxKDEPdp/
X401NMSuFg4QiJC713U2PlMoHVNizGCyvnL9qq9JwSzNUv7wYFNaEg46Jioxh95om3IRR6Y26Tbc
o7bzkhytbNLII266D6vd0U1clNstSZQshX5dKlAAEv5ITe52SI1iEMH0kfBH3K4PomTafnyiEr0m
sU5PICZcQGkbn6uXLLMyVLIjhoryx2jWQGCUcefd1CjUHO3NQdlhSq3fUU6uIWVXFt+mqzaV7eU2
wMpe0CsEqEknY4t1dReXGqS1nFtg4xTsDUboAKrZCiLbhE+s5LnTXVlLsp7hM4PTXwbm3lJwRs9p
4QmhzIUBVCR6VIPZaTWPwTKhEU6WG6U+8c7koVPXWELi+BLxMYufcTuSSZZbgYGJG2tj5EfTKVYH
a9u32VwFUHAUkYra+mdTYRfcDzzdVsaz0uIw7GCieyQL5FIuE4kXXrDCzOOgTyfBNYP9oatYSGRP
2D2atNAjTq8dpYgLEk1YPzVf2I4DFvpV29rt8CDN37H3O5cRlCYf8QjVm9GvJM//+UWit0HjpSnx
TEtpGydddzMRAc2ZfuzdxR+WsG4hixo7sxyvcQEzW3P9tddUhU/f7WDY9HJARjldTFg2sPUdiKyx
3GGONGNkwT5gZw40zUJlHcPGDpc0Xa8qtwZKk8gMYBr3r17Edw9WfoNmjmu3N0t2BlsqYSmbd7dW
yAHcskACrGsPGPTNMZ5jRIe5wQgx5DH/DrmXQWdU3obloWxYTvqd0Gwb6v4wUvFxWwcFTFFPRFjr
KlFlYtNdmma5DyiDtoLd8Tx+tOnLpoFeUmUTisN0hBzBYVIV9Cxj/gFrKYAP0wRyBucnCzUz69Nq
kJ4WoNMgTMVcLki8gIwEPeyJZBDs+O/12NgDM/Hq5EyZ0Bud4bXcqgBTiLi1A914ag0lROVVxzwN
HTb0YVFB2eaGhEBK/eV4lzoVaDzkgSrJFKuw9ZPrXnVzYjcX6rTbGfeA9rqNvaeZGLSw4LFX7+we
CN43Dak+7uvFMauLQ5nvkzhT6XS0LY/+8QovGNZ0HM4W0nrWt6qqyMs/8uCqOzGSMxSPA1Jv2Rxl
8NER2CNeqPIHpZ7seQww9EIxXyojNST3O2vzXuDQOEJezH9m68wB9HDI9iKypGPemhG2ty0oUujB
eC1M8DyK6xVLj3d0Lmye1ihndVYn189/3KgMhq8ZYSxh7vX2nZJ6I/+ly1Zm6bnarLpuBGpvgq8x
enqPbMHuQIMurxcXwvzWyWTgDjazYzTu4pwCLQsJhFN/Yjifu+Sxj7q0XdfKMfkAyHHolKJXG27h
8orGSuV04Dr2CCal1FfH0I85510CPtXYdPel763GUvw6oKpMLbraXg3Ow2/nUp33HFVQXez8AK/7
bHSfXrwFoWMbCVmzP+ql5cdHspybe0XAhkBdZigjDFJVLrXBj3JAdA8CIspiXNOcNCY9VGBcO9fG
nr/mKwf+BYM8cOeDmh3IdqzebOw0kgejAHr6xCVq6W7HaZZx9n06LE7UrM13kV9WS62B5IGBjGhF
iGrblzSKlhoSEZf8FgdR3Fr0DH6FNva4OnGcTniFcsnFuNtxxYeJdh9G3mJ8y8m6oGgLYvVHXqh8
/2WStZ0r+a+bNMkE7RV7fopecBJFVOJ3YdpeGx7eEG6kMj2Kvb8aydjBQpgsGzIrwi3DH9Ggzpcv
jdXoixFUNhYjQV14LGeFThAYOhkDyclYx7Mo0bxUiJGhhJ7RS2Er6CVGPXkf6JJdU8wTWYRpSYgv
VoOAVxQF7LSurTAKZXuafZkTi9IkmksMCPPExdvL0yuIw74vQV6GrHC/KH0DStI5PKHl+lBpX8Vl
nnUF2h67LMa9DRMrDiE8WT7dGCJLI4xNskq+A2ac+j5RHzDVWytitzBUDa4J7Reowyh1USnJies4
OOUJKTSPjuANv6hN+39ur3Krxjzo5B+vo+Y7yGWIjeGaE+J1LLbEawpKZ1/CF9NhCn4S5IoQ6KI+
1SnJ1k5OyELflZ2hhnwNatZVE5BSHsD6ZQRtTmxIKle/eVH8CUa71v3vSXu0XslyurYp/AEoQoli
xcHIircDXnurnxjDU54fYQ4dSKLu+GSUpZ+xn+HL7B7bKDn5CUG70zjALpDCI81eejLFJT7FsW9S
JpI8NunUutOv/xgonsJxzLjcYJQhK9q2JOTf7YTQkBUcZLbtQ2gwy4EZUnTTl/IIBLOAAbSfy4oN
TJhx1mYoCG9NddcbRlVLFpCXUV9c59tDGnDB+ouj2Sa24kCVO3Xw/hRnawbdxKYPzEXJo+yv7TmJ
qXnpdulsmsl9Ov2Uefa1a8bmQYS2O0p/kWV4WBQUeN1b2Ca35Is2MgeXpM5l83tqQ9Sz7rTQ0PPJ
24YWWAnqegvlOLxgyTCJceqBX88KTsOOpM46xfujogTPe6RILfhjPZJ/CZ2GYUQT3S9TCumuKdji
9MQZ5xhHxq745NQR6tMIpQQ149l96Mdr+gEQY6cvgZtbE1iTDCqi9CV5/Z3VoNTO6t7uM+rJrA63
N7aIqAYEMbGl/R/uA+2wFvqtSk1lenZybS03/ACnMU97qUKKW3bf7H46KipSLtXFjiao3mhsTGDR
ZgQpqre1G5j+UEVzWsRFg4bm92g/Lu9iBqhj2BCRnwylhT2ci7E0aux3HiXUibgW7Q+QbJmC+EpD
fRyBceaRrtgvllIBJoXsiFU3RMW0pKXBImBiYr6VgkCxiVvn9CO6OdC5DARAZnSLRfQhuZWusmFh
FE9ZoagmfYiDxovexVwxWunDoOxQO4963JhMEMLL7Wsk9xe6e26J9L8RKsRhpRzOg+nzaDE82MiJ
im9RnP1sBNyK9L5KjyHeuP8P3GvWOiqEgZ0oLHbv7VhK5YVgpFSRqlX/iLLpwXZZiCR60Vc64bnB
u9BwS25Zb+dOtbo7e0sVNRSAU3kTS3uVMUt3QrBywXioOPNd2VDwv5T3eVQj7Z+F3HVgun2Q+vXA
vJN9fOzG9X5f4OHKkCX+ULsv/dwir3lmBl93blf/VKoFdK5VAdZTFuwOIbtybrzC+t0sVZaiNq4Y
2xupqVEb1a5EagVoiXRtIoQhppA6xdQ6oZoFj4LHU9mqXP8Cfge0qI74978NGsSNJZFuboMGFMQL
HlclHHZHy1qnDTd9bHlPoBHf8xtczXXdjMzHt1n93u1WrMbxQ5jwzBdcE1htNRdU61jqCTBD08ak
bZDFSjCexPX4v7unPpsNiLBuizR1KH2u2mMP4T1QktslCz2vwF3GjxFxRfsayGOeMPBGMmdjeWD6
6BImYMRJx7il5+LKW85AmYhRUwttB1g7TDcOnCm0GQdbIaZFitGmJDbgl4oF7XZZYZY9b3kj5TcT
Q7pYGKdWzvrdmxKbWP56VDUASN8XYDZnzU+3wa+jo5VglZC+6G+5JsZAwhnxjVmQuevelhNlxzuW
7IZgNiwYhLWDf/r257yE6UipFuYF4zeRTN3OZJqGH6I4RHTUXhrXiaKplif+5o48kyJDHjt5xj+n
rPgAvQ9b+WO9dxNC7u730d0/JKo/MRXrnAakBf1L7dD7u3Qm0OE0DLkaslUqDYwhzZCbfRFZr77G
7Ij3Y4tekWYpzclKBCqoeLvbgfqrYQoWFhh+gCA+wBqNgM60ejSC0uXpkME324OLeQXvThhpTQ90
PpJv1IikDc+jMKAMhkQNh5tAafh/umhzO8f68U6zqiPf8gi59t/51lQkl3SlVIME70ZgX7BnA0W5
ACzuAo8KYzCOIiB/TqDIx/B6/qtpbkSprwL7Mvp9JLSHn8f2SZAhcOESOKAdCcWNF44GAqj879yu
PvmstJ3S0TrY/U6lwJlGEPfSP8QYnJgVHQAbqGSMG572k0Nz1vkUqQOoyuZUjSZnZ/xe93yRggh7
T4pr+9pTk6hH6pRVmJxRsAUcCP9vhQIS6BmJza9RsFFIx1Zuwz2XO8xPUgc50Q45lR7rw20VbHUK
w1teMcqLBWleRT2yG9HYdFTs42OH9hWTYm9GAC40iVzsT0VKWP+CVO92HT6BH88xHDTjO1yvHMQM
kRVu/N8Ikb6kzSOayXSZ7pRVZvlZaSKW/8E2s6Etu9Yn8uWx0tzg7VOmgblRkPtwCuYAGxxtT9B1
4KVb2yw8vT2fGCt5lBIA5Sn4fO1svE1zUiMXzqigRAiG7qn2I6VKXwCPBKVs4Sbevfo1kZNO7Vli
ioOXNjOczUM8XB+O94+N04uS3nTihEfVFKyGK42W2mU8JU4+g3yeUd5/Cl/g5o62jncblHS3Q06i
xK2mtZxP5CbWitDUkt9wumEb+QJFMvgXNpRwcg7Wp0vr4cIXWyWKQyiW4cJG1W1ny1RvoHZ0n8B8
jo7tB/rbGPVh2T3HCxYLj3fh/2H/94lLs398zFxoBHW4rVWAtaDh7mryCXI7mBLceZweLYsKxe8K
LXPjnOF532tz8ctj4eEzRArBemgGCsE2yId9WQH5Z0KiW6q4K1+4mTI3gscEBYmaY+sMrdS8e9MW
Mz4efs3Sf+lYwZrR/iFEtvXeEW84XXsg1aXX7fUYVHE1yHBdla/0Zea5G4Hrz57XvngPAQs42z3o
SezjoMun7ZnUGcXkL5a3V5Qrp5SUZdMonR2fl+NQSiw1Nr55u2SmN+272LBRYNcSarOhPqRCAH3h
WbxVLESCqf8+C2YqcMSd3r9OFkGROFzXdqmQh3z2LusqS2Qp5lflvps1GNAzpGDf47CCtwCT9uCv
c8Jj3iNEyO3qjfdEmF+QXv7W0ZUiviODITKQ7kEgZx83OKCA2wqOuiUP4Td+xg3OR0q4XNSfzM4Q
JkQYUaps92Y/5FjciKhCURL37sknI+rzQz1wUZrQY55NvCy/F3WtWKRzp4G0SqZwbKhu0Qz7lx51
F0FntE4575hV7aG2WRhm6bkFLTCOkpkfH4W487Uz1cHgsXZBT6drKdZ+BiOXIOWQQyjDIx+rImuQ
0CcESGiX6Y7Hdopm1G7lNT7G1xT9PsYRv0I8OfxVUmVtEcGeGJgDTkgZC4pzODkohswMDl1DbNyZ
3hPXfU1xkcbfrLpdh2Rw6Pilqnci+mbuStL7mUxCLGYEEulT1IHAg69s2dd5FbYRCioq42w/6aCE
kRNhNrYfnqQhjf3KzYeuYJBuMhuAOwZrFuZm1P7SigP4xucImlCR5c2rwemDjPNELo5nhxwQxE+N
6gLWrVs7fmvocDiW14T9K7ow8WkxklzdhDse3K1gr31e+2plGyq5qOCySm0nPUX4FnlUgEo9DdMq
hCmotDCqIqwKC7J96ucIJvcav/DwGz2yv3dVkc4fjAJESUMpZniJk/zvdidvFqmqdcO4TCOS9bm7
iIR6EahLjGbjYkJYe2IRmsX0oJuxieg2NSTb1xMwv06phN4xHtz1mc0xNGmlRm0sPHG66XxXKzhN
SZ/IiMLTt+aoHQ3pew1f17sKs7+7n0/YGv0Tp9No4UClZmrpv4RkPbTkTI+lCOewe1iq+6Z8DKeH
xjBrMtxPRYXbRAnJFLn7+bbDbtMtZZW7dqNdjyw/P7mluXxlS6jyp0jUkCX80RRTBl9tsdq9G+FQ
k8jRpjU0hLbcK3mQcyadmeRZJ++8QR2nlC8Q9cVBRvZmACGjtvrQJ4y2WtVueAKBPh9haLkhktUa
HSMbOa6JkSJT04GIC/zVst5YowTSW+tR1zKgdD++bBopAnnWVbHoBlFdz0BSYX3sxtrbhkxO8Asw
LxYWTk4m8ljdXGYXttcpPh3wXf/Nk9l63WY84ClUGIOGl0ymNkIu/LvWhFJCrxPWd5uhg9KLPOOW
6NG6w/XZfwsuxC0oE/ycpbC2+gPhb+FhWJkT3AHX7p3lY+DTzjly+CMo6Lm8J0LsBD1GGoZjwYkI
PWojx5jdMEf18U3x0uSw55xC4gY3To1Cuubv/fzmqIzwDVcgXRFICn7vyP+ecZ8iVPCPBYixE9bd
2F/aJgmdhDZIpwAR8/mUnhiuZ0S7Yd42O+o/UpaM9x8Nz3rqlWfrC8S7f/NwTCzgH/X3DtkPEr/F
UNMvvKopvOjWWNpQcVQmypuBXMKpsA14qpSy4AC18WFL4OjDeryiNBE2xBicpJefiohTHmapVuFd
2ZvMsp41o79rBOyhUPxISoLN7KE6eCPTrKQCckJLgwVkZa94zeJfwOFBCIs9bWxM8y1imFtAOgYs
kYatDOMm7Omvf/yvhyNdA9FJLVfNFEDa0aeug1g4+/Ww45+iDu86mLEE5qNVsoHvNBFyWyy/CM1p
Kp8diZ6JPQa7PBISxOfjyVKdCzHGtKjV8WITDXXtVjDo800c/Jj7aG4sCMSXzBjesvg+ShwC7ePk
oQIt5sYklZJlL6VQfblp+BqJGUDnRhcdJ6DecBzHJRuNyFPzBtEC54+nl/NmACJHlti0PdIYNQdK
Ym7MBfZTH7hhXQR0cOHmPdf2s2qNbl+hj/+bUsuW9FhwhCWME3CAAN9dUo9ZckZMKpINvCCP4EsD
XOm/wjo/9N3TtiUGm9jjx/z1R3GRUqOvnmWR0vN9X2oSOIpxewM+VIPonprK/2Kif5VLIh2g0/kR
fnVyK21DJa2WCJaPDA14FeY9YvAiN6FYSmAOlJNvhH+5ZtpRAjwkajuqUtyTv142Wyzqzen/S74K
l4kSuzIUZHg0SzAgt7yCGGcBZy0g66EDVqAPtXFG7BL6rSd4h9LGbZ8pMY8sMcy+bb4aeiP+L5xq
71MscVkCGMMQxJlHVre9ENtM6tFKgGY69/78VAkYK5vJKnSQNzV2SFGD5LYd/lvXZV0p3xyps1kI
O7bO9zhJLOi96H6WsdsHY/HiAyXMnaNbmDsOQscqfmlZ3pd5FBWqRVHfogxVjop2nYxlFMQqgHat
E8Mrz+JkHu/lesyzvV7DPAobX9Q6jnAkgwtES09eEIFohbBrweNrpvs874fNNXJ4Tj0xnnVqSYOW
ldWwdJJ60hKu2MO7xS5bWKTpR9t7lhZcwsjTFdN8L7f2CNgJr9TA4jz0irES0TuXWpV0snUTEyy1
/E8CNRCyVPJPOOcZ9XTNSlkLPC5uwCEHOT7+FlWxt6U2USgqub2x7zyhhiTGoS5tL4CMhoLmnAWY
enP80ywC8NkJGDuMmBmsOqyN1w4QkMg5AkIb+BGYs//GK66NuI/kkfwwDvdAJ9j6eeXS1jssKdAq
1qGITZKcURYotUU6NP/x2I0wtmHvpf+rx8adxFbyCc/7+E00JxJtJU9Pg3+s+nTPyAs2WHu+4+lS
GAOlLccfD2kch/siORibkseRnEwz5I47unTzfDIg5vbEv+eDWGwBG904MYmmvz7iVvnqwpYCvr0p
8mbZv1xQMheoeAOJkfOz/uoi/5E/XP57PgQkPLF0xvSE5AW3QMARcX1qdZFerokKym+phKorWzLl
0paWSUpUDTyebyI7axT9eCzc2ALmehvDAzPWQQEOg/l3hb8gJTGdVWQoc8BAQdaY3DSFq2VPFo5d
YcxrkTErrV72LNF6Uhf+RvQNj+n1U9PPGF75DIcqBWwis7q0ax+B/iclaIyofECIjJfav5yhRSQ5
3xghFqH9GdiQ6gSh9cLu4Qu9eR/7kNBtNtzMizOAUWIJsED7UYcXTBrxqkPDbj+0N+2ZU5ii8Ps6
SBrhgoqPewX7cc52gbh69EW9uy+6kkvZBZLviCvWvDPP95lw/CSgQBA8IHTr0X6ErxWCEB/B2XBW
y+InMRKckVoX3DG5VxZjuFuia0KhviRwTAtLHs82/mXebUQZC3UL8dL3AnfClUI9e4o2yBMPFa75
ywowfSv9g1hw19HowVt0tQR858NcH5s/4UAZwnnJBkfioXOn48/5YogVZxZJP6EScj1EjlR3gS4w
YRi8Ze4BVV810MWb2fGlE4x+o1YspSnqcURV0sR8qmLiasbTYIHrdXE3KzfgfzFz+tgL9cP1z46d
qwzp4+3LzhAe7hV2evgqPpuwFFVkX+SiHifwJSwLUZZ8seKfblUJqMj3oDpfrisi5bKHihGAWNzc
0jOef7JSbAXycSC3X8fAKPGdxtbNVIYvZpbcmh7K4xXwEzGaVwRg0qL9H/CyhLHOxPUIfCxMl+W6
vTfNzLhRGIe31wxPKMxNjSzeArOK1AvRr0+ULmyruVlW0++QDYI1YjdisP41CCbkHfpHiMojwwb8
AcGEAOzAMRWI4HCEdTnWefOo2XDkqJMkoDhf0z/Oe4jRedH1Fmuz/7TaWUQQ8iBOlrfIPg4cO4DB
5PkPHGs+6cNP0djeyxvggiWh5KHdPWny/tnj6MgnfKV2Wp0moMu5nBQzsDs9/F+oZcrOFzyQlObd
mNf36BJD5iBdsJ9hxiCZBjgOpBdlB3pE4W3Z1s+iZdg91t7/UYUeOUjiotBTSZRpSCVqY+zjG3FD
+6u8b9DpR9gMM++RyS09PX12FTAaEg1D+LuIy7pFZiGbIcSgyt3Xjv+56FMuU5b8SgKeWpvCjq8D
7vT5RyWwHsQpf5O+hREbu4nESW5n7FMrNbLBsnV2ir1nxqgVLQhVEcuvP99bYxWAeZC86JWKCFxz
JdNtqA6Tuup5cTc9iJcYH20yC1zslCr5ZLGAX6Qm9lgluX504tMyg7ySmLBM4cU7g8gRTqbyfVvR
dddEkjz9i3IC/rmFaXI1utj/xb8YYFYXA9d8nN+IgMvI/zRqDY0sbVNnVEeF/kug+jXz1aD4tc5K
n0Z4TFJorxPw06RqL5sgiL5EraovQWCTjJcfKEB9dZYrunL1peuy92RQTndQik81g37r+Mugo2NA
OZub3/YYywOZ+hG5STsa/nIFfvmji0JoZu0ZaI/9yJmqHRukR/nw3t6hTC2mNAuxMIEmGYEIO8YI
lig+ShH64ZTOzzm4Wzl69vB4qSnJwqoYOEg4YJmUTBsV2aZv1S4eGQAUiqXEMYV3HFSuaaigYHMd
Ue6DMUAotqQ9yJw2tHsc5ITpKVf0xwArsoczkGIjh27MkIXWCPjANWebn08my/X1byXlq0nPE3ml
kLTcRdXlwU3QdglSwn5OFdyhdUnDso7wUpL3Kl3XnTfVGWgr16X3ApgV+2W4+T66jiyPPED+MOS+
4jaY7f7EPRF7U1NwaaYb2jk59sw5+rdmXN9TLHteisU9aDkHoEJykVb1X8pIPAUQcaZt2nt1HkGY
REQISnx4DuLl4K4uvn1lV0rqIzgOLDkEdEC/Xw0FjB4C/WxAOhjbYkcgGgys08ShJ4MStOjRmuvq
fiq6dYRwSESacWdazytbSlyXuE1iNlBF/20uQvknBzJok92bW3bMMDOF8Hcif6x/vRJ65vPvEkAz
dN6Qo5CbMBHwXAE97A+eGNt6jjt/AmFMV3ifnNCVTUT1T/wDd0GOr92JRv19dnDWrfX5wyS/XJ7R
inxsSGLvynf3rLawsVgNLBwUvi+js/znFKpYqd8bpW5xGo/7w3io0F2l/OBiHeTz/bGZCHqcLZYS
wMEb9cPomNc6ZAXwz5iFNyU768ey7jNBnTMVJ3qHRrWO8XxD6PuD1u/+c7rs1PU6fjaYaUYaq5rg
tA6zvxCDRXkV08oiYE2zY/Unx/Iocp1Ib2g6zBISW967UFoBE3M73NYUyLKY7cVCKl/mtaS7Lf43
HfMVIL4tlGF1CcaB3ewFZDluQ8ybR8xOX/4TxGsHnpbX68tBkCRPrBkHPskTDVhMydc+8MJkJLjb
z3YKtU3f2Lf1u3j37cwOk8J2YdQ+SE7XWvRuz8rFysNPhv7aMG5i2scv3gtGWjzxgtzEZpFRAoJl
xw4Z+IU3LHjEccRIBxT8ykrwbAxLrcQGApuwSPTiXneeF/viU7+DZMylk35Rl40Wf87RAjc/KUrd
E5hi+kcR6UVnP80AKYYB1qTJSJtWvIBs3HyLWrGDFpZTQOpKzwd1xFpveXOMaa8lV0nSC0se5ygB
EwrOANbsfkNaytkouZT8KVYxJwLGMtGrBc+gcytoXlfAfCWhvHgEffyt5xOkw+IN3AFxDMbF6ASK
wer0Jwip8TE1Yf/2sT2BJrYK3wUaph3gmWpppq2QRuayG1On5rhXuT4nr3hdvp5+A7+OMwOW5Q3+
fuRYdWuML2L1P47kc4ugsrABvOWktorI3Oll2R3b2hmIXWy9Xnto/XrAhp92UFf/z6GrzugSewXQ
i8uqvsVCnn2FRP+0oEYVh0PdwvixVp7V/zDd6jagtSUrIfwFxI90JwxuE/RR8OmoQEcw4F3eXifL
Z7qnqmY7diAly2bOW4vn2D55e7lSJQjtpWPJLDNq9pfDPnG4vcn9K00nh3S22KgImOmt7hvkjG9Z
10hp7zijgNbeqDKCHbWoqTx1iEh3Nxz7vw+q3msp4H/z5JtsFIcDzj28EFVaz2SaW4U6hi3IcQmc
UhwsmN4CjFHxpCXu/S5i4Jwr4ZTAufKbRtOMmz0i0IKOzRmITgBmWyimpX7Y7vyfGCqkHJgfGZEv
n0W++aCS9P9vwi8xgZTnlWwXVobseBnK2RMDDmL3Ej2D+/z3nzhZR/57HKjzuR4la2A+Kr366xzy
xFVuTrvlDqrohIG34gNdQfFX1UPuwJ+AVBhFKfU19CH+MRB+huNdVPIqQOmstZ4xXfNbm+F24Dlw
ABY8UJmdXVDZVfEKvpgRvsv8BqiLzaGNgLZEcdWREYppM40+GB/ZYCwwekuHtI5u1qu4Mttij8um
I3iS4ht6wbDYX/oPWOLS7p/4FLM5jRluvV6sECAND68XQIW8Ji6FubT8mpp4BNZge+XqulJHYT8k
HNJkD9Jioq5Vfgwzr+9JYt5AgS9wQ9fuKaaICuJH68T41RVbKYTpnTpC35dREjXntGlWFdGsVz7y
AevitU1W/vEcRxoC4PHJ3z9RTpFq47/YtI7CaVP6bY5g9vCUPG7D+sGK+pNUEuJO0+IEgIhV60Lh
DiXi7u2WKaJfeUAMkIUO1Q5TTNvd6P6ftFqw4zl0l89Ph76H76jTjYUlaz2dcwXI+/acbFP15a17
ees8C4jiMjnLK/vX54jDOB4T/ZRzCfW9/FtStdty4BbSy9a7XsB/OECOREIieW0N3X+BJXe3TCEC
C/mNzo0t4d7ELn87G83204W46Fn0KztNdEmUo91JMmd1ziEqZUmsW2cqW16S/8QgdiVc97ctmI7k
MKSsLyPUJoGOB2Wroj7TIsCWaLMO7VPm/AlSLjJ+6GiUAwrUovOC2eWL1Mvi7dZ+7gGZECBLzhG4
YJcGNwA3vwuD3v8h00PrwK0LZKiirF1SvnXUnohlnG9XoAobUCxr/pUCqZ1EWS4fAUeO7R21ZW8W
Hg6L63xwc1L2L8e+VpDqgalfxVcJA/dFjamzu9OKdoTpdbQLeiJoP13WWfwBBIywRKGArWb7GqhP
wvtxUWrn3oyFTYEhJ+yCbneb/BG+eEFDu466KjH80z7SKRmC+6gDLg/NynR1rCnCYFqULy0LChoa
bGl1VOetrLa6QeJTkKTOUwav+aY4p3Vg7yVMvsbcc/PpOQmjkTFQFI2czuidX+sag+nuOqLZzoxw
EUI2Iib7jkTm04LKvYlYTWBWW+AHe1c5CPiZPx5tWRkuchD7B6kKr6ESBvtkk/otETrSXXHr6XGQ
h3II6IpUIntVx2x3E3fMuNXz/7KNOLBPAahWzhhEQtWfF9tJ7Se295emHKmRX31cv2rbp8oBwYdp
9irf4V2W0yg9jbpCHZnWDuYsmFYexFml+xFBXVvZ7maj8VDWIMaodd/Ki2y4WLKtdfj9XIjO39Ew
Aa6dEf0Qm4TUzT0P/OLBSDJlIw6nGlHQ7RZViddkWXY9YHhdz5PgLw/sPJ0k1XvpjdklKUbsZDqu
h3jzyS7iEJs2Es3JtWa7uvKbTawnT6Z8uaPDwgI0NOv2naaBVGyRKf6CWEw6Py8KRs1uV1TH32Yv
+yql00Hb26nyJ87oM1nh1x7Azd9OIBGmx9s1XFUkOOCzOI0mVUSQJ8J1074SgmJhTQqqLxHnm+eS
ciHShuitz2U4R9YAA2JVLvLkQ1+jR+MWwD/JCu6oyxZRZwOwN7x1WjOSkVODpl96/2MjtLg6utQl
+z9GHbasR+nVIXBcIrXcj6naNXU5xeLJ5ARd4Z4bCOHzJtwATzesLksQgENtdRDDTeGVjJ+7P5O3
wGc8S1PfmetACXNdk1NAd2WdU/OzdHhBTdODBU8Mfh3FQiUKR4noWrngJ8/X/HjT7dTAdS04XlP5
RiZfgM6vkKEO6qcOpnz7n/9CEct45faIDF+Nu5t1LgC9gSbww6v0eJbrtYW31JsRBLFKK55fCdbI
L2thD4NF3KQc2Q1u4LqolyEZrUSYhQ+qUymemKkGejm4lSOuxVrnvEnT27AHZpyLdywtj/Dd8Pxe
PnfnzSo0rU5ky0QoxyDveaIgecBbf+IzKOYBZuRrcxSYUmvJEaaK09F/kefOrHIXOtPKFUcPq49T
4EofHgca7JHCiLupT0+7+1KgEspyhFB7rQfBDYdi1Roe+8OHrUQFGcD0vk0bMcP0+xArN8INlIYe
KsoDogjGq/B9SHKHqwCis6PTyDHYsReKo7zR2+v7J5/C1qwHvq9CLPeq6G5p5eeSz1q6rPcjsT0Y
JomW8iW19QhEN2gqHaA8OE0RiVGVge1FTYqhwOsMc/iufGdPoREHSWF+ZQiiWG/Ju12H6hpkAUf7
DI4zTLmUhMg4TcslOdTPnx25q4Dy2ryEXJk7j2LIlLjlNoEfGrPJYLTdHXXmfMapm6VQWw/bvk6D
zf2SQ4l30WvBvCU9F1wywHnk/amr/HkOwEJBB+w2lt7SKJCv2nUGcsG27LQsobErQxi+BvYq5Yx3
wvMdwYADarmrC1BeHWLb4oaDbkDOw+bkRA//t2pHJIZYjkR6AS8nR/Gy4SZH6VR7QfWH+IpbwTnd
zP2IyUN2x5WF0qNy8RejNGZthLfb2VWT/7e4vY/tyU3E0iomt7h32vOs+Sun7ibVsIz+CpynEtET
0801lf0sqdFY1e0M5dUHzTlkJfpBZf1PjlonZDfVK7UNFlm3YgVce4CgeKaa8qsEvb4f8G/d3AIo
wB/rhn3D2VjYXVZJ3ZWuzMEbWIihSAr+UbwkDJZzNikt1OoChTTSh6vxpS7nYrPV42z76QAnItN2
6qP+MDpJcql0w7buj64OH1EFvZl2ENsycgBi7hz+Yq2uIotQWu1dFYzVleWBSpwuISKXqL0rZWJ2
gwn4DbeJW9BMhr5+jdus7OdPioY7Y47P8Bkrt9pvhumFyEMt2gPY/338QQwSGvZaEZHJYaoofqqd
kwjyjjJCbgTkKZ+rplghwM8gwsuoM+rBifAHHMr+/unmmoTi4PmPxqiL29uTyz3OeZVk95gAw8T0
9R7c1VbeNRqrJ1MBXOgKWzfxAsIUgiJyXwaTLG6ZPH0mIaAtS4hfhj5d6wra4WvROUGF4WZlld9/
ojl40vvTI1n497hM/GbELlVVClw6UJHWy0QN2fKpXlsGSG0wBFj2zVYPGkDfco91PNf+qmvlSxs/
pn2caSK/XtDUFKJKUB/AY6SC9MUDdNu7cUgIab4BAtFiFXSl8TG1Ew+x+RZ9sioUXXrxJ1lnpYPI
FuHAbuKW6BVCxmsXcU0oWmGfxvmkd9lTlnLemYCStt809S4GP91/ndpkGnc8qmqls3oveo9aq2/u
B77Bzj+WWGIkk7Chg7DeGpe3SV9CXK3V7iLSar+lwYiWtz8iyxoTFX+PDPPGJQPAYj64ZlhyktTM
9b8T8V9zc4oSXu3aC/X+gMU4agIB9YjJIF2uyg5JSClChoo/myMaSBjvFctDFGMhCNJfZLLp9cPQ
LQP0rwdsf4G97WHuLoa843h46x1l9Yx2NWtbJJO+eD6/CR/5KNFMh+sR9Q3uK8W6z3e+B3DJSE21
JXmezhKAXwAHjsKWhqjm9138PuzaujghiqpSe0SkVgDgpwBqZsfLUQD4AkcGKJUN0yRj7aytHeeu
+JNJJmiklI7+Wh0Oi8/5y8L75OIcs2LEvvmTxFs+z7r8tq3pFTSqYbP/meAJQ9MgTtGdGVpN0pwW
SpYWxcioiQQxN30hl9XkPOMsYz7QniSt7elhnfAi4LDkvRMK0FthDzGyxOMhCE0YZsg4smPJZXvj
bf4xc3xK1G3zrIpisJiBOcttroRp9SVOQORZR2AxEWmOITj6pxHBVbYEIXsCzAsGCn8hUe69Ld9c
GixBUdm8pzlKma1sjDLA39t6xwqKopFxwnUX+v3Kt/rRJkOCuEcoNFGWD+1uJobH6t4vTZYsToAi
jK0bmGv7aQtaRefsZHbhNmcPK9Ie9QUS84IlJCsBj5L6+NQghTzyJ56JZEMC7vR7kcciV091vkST
6gP8g7AkTKkZddg1yfO7aoXwypSYG6WV+/mErQkcWuxMXRD8hOqVz6RVvATb21x21Sm+074N/Fi6
oS+18SMmwbcVTxIjSymqnSUKp0V4JDrRsKh5DReRTAMbEhW0doGwgJJSyXKd6AdojKxO2wwO0HEJ
93tKaevaJOF42qe/1qV/j7OY8loYY+4pLth7hnqxVszsuSpoZVmMTl1uTfUYYjUDsrs9VZh9blZI
00//uqJ+IMAwm28QWtc+EZTyD8O8Np6VulIpUx+VPRBeP+bL+OmjTnjGa1NQ1Psoo9CRSt3Klt+v
7x+tdDhA6f2XAJ9SxQwmD6UPn6txweAVi/X+3+GwzeI4ZOIxBTwFCk4uUbQR9zS7oKQv20Np6FEj
n8qrsLEQkxAY16jW2CYLjRfb/ax5QvxBVY+JqRVWyuah6+mvZH2KEOAR5ewSMWMY3T1k1oVCUoQN
G0ofDyCFldnkQFGLYBylo5k28pZpVgw6G2AvYBzNO3rg0WnksESwT2b2Dv4pVeXvTQXeslHyCQ89
+amIi858uzn8LnKT8BkbrIvn/CB1s5GijyzKKwxUsB0InaW2jPldR/wbT3dqg+Pa1QpfuMaKSQod
HIArQP1zVkBISiIuK7xb8A63mPN6K3wa/qPfhR/RemI2ELkrExbf6iu8XTC82ltNsmDkyfXN73Ic
2kBs5Q3O49k1aMI99e48wmKw9DEYFHHUTo4N5WZs8MKdqQXV9xgJ0Ma9ltrSa9cRXQGo8MY/SDiz
EYJSqT/V9rvTg2xLJZ+8JT8zc8ysJr08qfbHDW/+0Z0XtIIMN7zIux7Owm9em56vaNviiPfjzut7
n/yV5D4yspiRvgL3cb+zeGT9Ph2Vefg1BNGDes1cvi6L5K/+uN22qB1sggyRyvc1/1Xqr4cs3iZo
wNzm2uf+7YtHvGzWlv5EIPxXGeYwyDo0YRw1KWkCDruMxq6FZDmIxYFHG4kqTVw+tBI61mMjfm0L
ieiBdlbpRmljy9WAUrdBNrxdXVYGqF803lfmHH/KdBQcoITbFXzSckI8oEYi+ZDVqKyEGnPVqMnt
282Imae1+zxeNR1SoDqROWhYSBh3I4A2cqehpBGS17xZM/ZEBRAlZx48kCCjQfwlEy47idTfL0Cu
33KsQtityBhghvdR0XiPobhij7UHU8W5Lcs4uSQSwgoYAM8zXpKjt3oaRivTBw==
`protect end_protected
