��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	���v�T��_��\�F���&Q�?,�xf���4v�zm^7�o?�π���{�D�t��^�aMH��b��DJ���N���&��	C�Li�|^ce�����itֵ>.&~�J�
m�~v<`��̾��l���K�{5�qZ�[���8�g�`�� ��n:tYK�0<D,؂B`�����o�I�a} ��Q�V|x��~a
��R���M��6��"�2��3��$�U��&�4�\��(.�ڶ>��?�@�2�mA6���3_�z�wC��+`}�l�8W&׸l���9&>��6%��e_MD8�ː9ѡ�2�"��M�'MK	,r,-5i҉�o�Ham��`�w3$�O0�?#$��>�υ�uN�j���A~���H�E)!�*��!�ݗ�/��Z��}�L4v��%�I��W
R
�Z��}B�X�Z p�ڤ���st;��7��7�@�|(N�!�E�� �8�e��TH{�m�l>��A������"���r?������!@���B�g�f��Lj��t��UB�a)�Ͻ-nj2��2Ȩ6�����iUG���Nߢ�2�D@�Ѳ4`���Y�)�.E+^_Z�de,/0ȟ��i����%�ܶkp`_Ҳ�n���h� ������kQ��)�釚�-�D��Lc�0�U������s��[��P�A!_�}�u����C1�'Z�.��	0o@��orؿl=P�0
< ��H�� �-!Py�&�A��^*1RMRUzv�\V@d�R�+��j7j�Զ�s��(j� ǫ+|�[�au˚����-��4iC)�4̹K1�G��6��Zʥ���t��-���9\� ���vI��T�[�S`��md�9G��Z�/n��&��P���+����6;�a��r��}��S8�]��:�~��F=��C�h�3lk���8��-�3�-�����IBY��]|ށc���slĊ@��RgaӃ�$P)�Ln�eB�t���*!�#/��.�z#�qכ�g��Tt��D��&����{'h�S��-	z�L׽��G�@�_&��bV�]���![*��o�0[�{�gy��lG<�(k�� �t +��^D����[�2zfD�f �����Zu������21�`+Jq�����ע8y1����[����}@)=����!�q@�O`�{ދ�AI���ߞ_�ƭ~AC&���nE�l��cr(�2$7�n}k)8��v�_zC�ކP�n���4O��ͼ!5rN�d����T�`�y	wW*Н���#����*�&�4�?�t�����dC}�kn
Q����6��ki�������on���}9�ªs����\&]�����CCp���pa�#���SM�~�U���]|�����@L�p� Āt���H��N*�]Xҫy'�Ph.q`�����Ɓ���4��y���L�B2\���C�mT!s�Ԣ�͆s��(wLQ�8g��@.v�8r�&N���N�D��ܴ��f��u]�KQ"�j� r�v۲����fȋ�L�5��?�u�݆r,�\^"���Q�j��`:�Y��}���DؖkA<�^`B��;�ۇ��(eZy�S�F�����˞\�F��Z�=46��2_���L;����p���l�E�+4K�ݴ�i�o~�8e�w���
��'|�o].�&<O���e�i*o�eS}�]�o���c��zi�[�b/o�K��"o�s�p��΋�P��no�.%��ڠ ����7r^�Qf���"��t���Z���?v2�����]y'��&\f�D�^�E�����}xdԔ��sבAdU1�{�]+�{���{
b�66؛�t��pHz�vc��[�̅�ϪR���ٜ	�1F�.ab��7	Kó�
��H����!<��T��m�?�
����Z�Y�#[Եu@��C�����cF�PK��k27s�&��~���J%`�V�<��&z�U�"4���!0�ƺ���
؆{ڈ�L��h��<ړ�)�N�&�}�5�|���q�\3-A��1�$�_.��D�) �fWsd��/�S�ƕ��$"���P�u�Np
g �N�.�Q� i�7� �#nc����{�UC[�CX�pK?�7��0C@���I�R���4?4v.�!jp��ѓJ��:��~��J"O�!�+�/.���Pʰ;Ќ,�X}�)ڷ�5���زC�c:Ri�(�+�Tp{L��2Tbx2�3�Սcϓ�_�j$��%���tq\��bwes��6ε�Gw��c�[�˟��Ht�z=��z$}�ț�E�ko��ᏱP��"ںG�C�'H�ԉy����LM����A��mMW�����l�+�������0��ǰḢ\Ŵ�Η3�QßkB�X�3/���s6B)�D>��+{�Ȩs"e7g�����^�P�����|���Sh�����ôAI(q�ƭ�gdO�n�!��d���M�M�+�ˎ_%1Zn˂���"B`Ps}��$^�<W��೺^����{�q�uk٪��[&���n��B9^Ӝ����X�?�j�֟)~ls�AAi�\�
��5K�	�p����}��]��p�%ĵ�JE{b��k�wn�����qG�Ӝ%�z܋��7��FIfI���n���yp�<�@�:���	w�i���VT�4���Ė�t��T�C���eȊ5A��@r!�~���H�%Ҽ�"�֣v��� ;�
X:�i����5}�YV�����E>�ʭdB�~� U����z[iė_��tE������(=����2����Ɛ�&;1�-�E<��������r;C������퇠���Y)�fG�ITXЧ؃i2�W=��7��_2+��>�f��K@⩀_���I��wi���S��O��!`a�����K"�K���|���Б�
�tF/��Y���^*�<�P�V�5������
5�n�	��t�?��6�:�����J;W�� �'����t��&.+�D����Q��uA>�a�j\�1�5����C=�zp+��t�ȭ�	b�k�R�g���<��A~9��c�a����a����rX6nX��F ��ҺY�L��r���ⱕ!�.��{b� t��ը�4f_�"�(y5�ہ^>
�����d��NQ^VTY#p[|B9�V%���:%fV�a�6����_�XYш+��^���!��e-��U5�T�uՌ�6�$?�(�R�����y��It�$���p� �i����Z8ѱN��,p�rN�`�**�&l,�g���RY����k߹�M�2;eg�b�ٷ\������]A�Љ7�Z��|�;A�(�`뢄3��{N�꽺�*ҝ(R���
���C:��3�P��z
����B0�~J�]57���P#.�d��>�{�0�����rX4�Z�[��6;6q�JO��-�x���i�Y���2�v]g�f������(:�b�^`�tD��a�)�9]Ƕ��t�U7�˘Q���]���k,0��&R�f��^U~{��>�����=F8=e�QtQ/�d}�������!�⡠��a�!F�ő�Ƹk���6{�\t�	�n�o��q�+�������jm�`6�Pt�<,3������ G	A7,���DUZzc0��B)cN�����+)˹ƶ��\����>�=�}6<��yҴה�a�"Rt�D$Pj+x�ɖdz����KP+�̺��@F�M�]��@a��L��w��3~���駎ĘLW"x?Ox@9�|�3.��~��*,���\�S��q@;�d����(����S7��K�U��$xg	�[��B���������Pw l���tsy�g�$������¾?�aq?�b���Ұ.GD�J4P"�w��/���	Y��4X�#ݻ�(��L�[b�6~]��H��ڢA�6����4�/q�9���M�S���� �Y:�DT�`�+�<���:��E�q8l��S��9G��Md	�Ut�*�p�M��Kd��M�e�M��.� ��<�i7�	�9C�>�|����B.�]e	��m{d���Ӵ�[�������U����<'�cek*߭�G��ڳ���ʋ2�6�������w�,�/py�3�!n/���|ð�Ζ}bfK?p��z�9��S��A���-Jon��¥іfx8����ր1����,�J\7Ȫz�T�n {,N�����,���l���x���m�P����,Th�?����z��mj#�2��T�<H9���q��uI|�����.!,��kyb��23�h�i��R�\��OuCJK�,�E*�6�ɑ���2 �0��F��B�"f
`,bN�	��>/�NB� A��y���DIߧp
B�d<�+}��7n`��N��(V�La������x�+�q���7l� ��Onٿ )kW�.N}n4�T�#B�.Ŷ���,\��_�Kv��cξ��MV�p��ͤ�~�#�J��F���������$ݎoh����=�I޶Z�����I��P@Z�>^ƫ#�I����r4N����I�P<����S�XDp�����7ڟ�R��{�U�>� A3p ��5%e+�ہP/����
�huDQ�ظ��65VO�6��:^+=i��eЌ��=�j�3�ƌdPF���؄��!��Ma�{�?���� `�O�e���L�j���LJ#\�����S�ң�G��������p�:�j�+�G~(�8:�I�]�{�r��0�cJ�u�+'�2��,U��Ѫ/���D0�뽾��*Hw��"y~6��pn�����V�<AN�p��2pq�*B�Ԫ�Q�^J5,DEs��w��/�BdlAB(��E�}R�N���A�X�#=|N� -��es�wf��y�d�H醰"��G�j痋�o6J�M~\��4�@0�/�e�S���Ka�V�#�q��\k~u�Wfj��(��8�x��8�W�Y	�C|���#$�n�yS[��!H�3q$k�w��6�����^�5P?���p
�c���Z������E�FP��H ����z�-����s��ʕǱ�!izi��,>�^��^�D0!m���[�عu�	-h�<��MC8�r
{�4(�E�Ⱦ��U�љ)T�p�RC�l�~��IQ�8+���j3q��WW(��&A'�d���e˨h��:H�'��>�x�7�����/�k|'3|Gi�Z]Xʘ���5<{{��K�Q)�3��r
��Me��,�d<U�����	b[��G;n��%7M^E�QK�v�Ӏ���1�*��z%��)��`ԡT�J揷��Ӂ��l?���G�i�����e���ϥpLя	� $�Ş�CL�B�����p4��:��r6V��W|�BlJ�D�h���ĺf�&���	(�qt�k�b�P4?�>Φk�*�}�;՝�:�-���e�"s�K$�y2��?���*��,�ly�C�b?C6_nCL$�?/�Ű"�3�L���:SÉ��P�ַ�B5�T ':g3�^9��u��H#Td���]�t&��Y
\��u��U���D"��6�Zb{*PU9^D�������u5�~�L�r+J#t$f��k�6D���Z�1�)���H��qQ�~,X��ɓa6=Ǒ$g��k=���BZ��"�`,�hsL��im|��+M��J��;���w���y��^Z$��_Js'e5�}�x�ado�R�fd�)�*�Z���2->vf{�,= ����+�|�[�!
Vr$:���>6̑��pQe�A�֪`�p�Nʌ� ��-۩��#�d���,{�%#^��B���Q�A�ϛ`���\E��l J0�[k|�Vl��:e�JK&���xmR�' p�u04����>@��踔�G��k#9���pr7��o���C�o����{c�m��j��;	�r����
3�X����N�(�nO��ӷ���gE����? ��Og�����	aP.�҅�������n0̩}o�9�Ŭ�,��t��K���ԅ��	�1OTA'k%�Vd"LTSOF���K�嶭�J�eh�
X��z�"އ��1�"2i#��-���ɘ2�#)PW�w�}�K_}�?�JVo����ҭ��eܝ10�������1'�9n�$	��#��	�qkM�܁����@8�rɍK����o�[�Ft���u���,<�����L-0�Q_PRy=�ͱn���2�	yx%�r>� �K+�#W�0�,���%8����tr���]������ް���8��j�Q�H5A�����~#��:���j���O�K}vj�;{�v0k��>�0���9X���펼ߪ���e)�\vs��9��bT��/٦��!��L�����x�~���p�Pr��5��t��n���V8��8������=e���l�z��R�_�,6��/��Mu�7�)��ۮЇM�.=ᘕ+*7L���6b�7����R���ʲ�5�O;�7:j��T������)Γ\�Ĉ(Not}�f��4�~R+��^�?A�����+	v]5����$�,�"� z�^j�E3zM0G��9���� ۠F�tևteuQ@��L_'�^�di�C�Wy�9xf�Ď*�����(�F�]e���S���jC3�L�=Ӿ��0���
�`��w"p� c
�=
�1��ѸQ�����GE�چ퍅D��L�r{Pog�p��W��y\��Mǁ�T���OR�+�9b� ,���|���\?�6k���ʐ�=�Z{;;f��nU�;3!�y��ē�&6O����'�`ϘzP]duG�=��qT����E�ԏ��*=Y�+��@n��I���&�:e�gRN�I5�����#VV��=}���9�B�f� ���_}̃����-:��$�ts�'GY�o,2��L�_Ӊab;9T:�l	Z�4}�]�:j�Kr�-�H�����o�o��4��ʎo����V�"����}?u��H�h��=1�z�`^eF	��j����:^���m5���W��x)M�	"I��{e_���Q�Z���}�d���ߩeh�L�*]�1|�c:�07�q�Al!���8Yѳ�C����I�E���'�m�����9�+O&uB�弛�L�h�C/E\T�B�b�q��2f�1�sbo�P�X���j����)vy��#t�9(E�|s�[^����ʵ�����}c�+R�5�ޣ�g�z�fӦ�ޫ�:��0M�V�4����4'۽ؚocp=�y>��t�#��S�m�{A��`53ۏ��,��0�`�.K
ӗ��K&�s�7�b4b�!�5D��e���8�����/�>^�z��ӷ#C��>�l4?��S�͚O�z�����^\e�<Nפ���t#BT��e:~��t�V<�B���U�S�>*D���1���9K�nÂ٠���u�N�����c��zJ�:���5_�%�Oj���51v`);�o���JN�f_�9����-!��������#C�����}!q)|�u,� �2����[������#��6�\���h�K{��tI��w��U�je_G�~\V�&34i��0��ҏ��e�gνɹ�V�- �E6�HU�C?�K��M�C|��nB�.��]�1���t��T�*r(���F��Ics����fT53͞?�2���`Y*�m�cv��<',�-\�{�3�v0,�+�+���}dw/]��-�/������ނ �ߝ�߂����������~1^~��Ty�᷅+��0^�jxu�����&�y�L5��J�$�65�]>��xS�X@���J�{�Au�w�m�lŨ:�H�d�M� ��&�/��9mH���C����	n��4Ӿ��YM�ŧەa��ig|~�n�}ݰG.�y�WQ&gE�z#�G_��y�:�z����֘�L%��+Ip�@�x��C��!)�aQ���c�����ַ�V���T���9˝�>MO4�Nr%��PG��������Ɋ��r�.N�Kn[U������4pR�6aq�X!v�=I�q��)��C��R*�L���S��1��՛�o�qM��������+0f��6/�L�>�:y��׆�B�s�z����u���Pz�7�i�(X"��vTI)S�vO��~��e���b�!*�#�f'��c(Ե]��R���{�I1WR��?�;�7���zy/O����u��%��2�����BIإ����{C�y) $S���c �ܝV�<�8q��2H�R���q��c��O�C�)��/f:5h��>�F�$���ǂ���允T[��sM�0[��Ʋɲ�9M6���=(?g6	����X��T�z��2�"c��E�cd���`�ϋ9,Z���N��Y�����8.6��XB�4�9���*^x����e������Y��w��C�6p~�\��-sQ0&TFm�H(�\f��)�X �
ĳ�Nk��2_@�:�(#uŭӕ�8�p���"��U�w=�q�~c��+яz(�󋈐�M���^��~X�r�	&&`�=	T�X4�v7�<�i�wW�������s�cdf������?%�'!_0{x��
"�7����v��	���\�~��B4��=m�-r�%+z�y[��[͘��y\z6�m2�xF� J�`h;F$T�Θ��6egi��o)U�[g[E�XV�LoD�-�К���zI
Fk�{�ӵ�g�PsЌ�q������}U:�B�92q��â3��g��B���6:2��>����nO��2*m���9jd�3/s��Yy����.tG������Qc��a�BZ�*x��q�pC���PN�#���"=���ż"N�P#S���y�