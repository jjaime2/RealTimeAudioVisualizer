��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊��Nwk-M�X�����al���A�[.�Vf(�{i�b�1��A������S�×�`iG����aD��Ɇp�2�"�;���d�����b���=����X�}Yާ7֠�A0��Wlr?X(�����}<�*��G�5}#u!|�f�I��>u�s�N�f�(er��d�rS���V���""m�A�|���� ��v�����P��r�]Q�;lk�������H�4O�iw:&- Ua�~�o�(�0�"�d�E�wա_[\҄t��)�c	ܘ]]H�Z鑄��̪����I�-��E�s]��=��������kD����3%^8�Q�~����e�!�Z�q"_���J�Tv����c�?KW�c��+��Uq'I+g�!�����-:��|�(5�����o�TH�n����	�DE�R.q�`�b���)�����>j���e�/���_���/�Lo��J�|o�!�N�چ\��v�/�#��=���ϕf��Q�n���n�SS{�)}[_��t�\+S_��ӭ_E}]6�1T%aZ~f�+�j�	����⏛��fb�����Xuh��<���o굇tЇ�7�#��Sؗ�b��C�����D%���3��"i�dif��$	p6!��%����_��YʂZ�� tw����ө�itܱwH�!����P��R�;A������i��🩥:X�=%�Xzȴ��'>��|�Fš+��lb���a�� ]�� 1���Z��qޝ�>����`�z�b�;�8�f���*�%tK�UπC]eֹ�A�f
�?�r|�:&���V꧷��1%������F櫉Dz�#V��y���x�e�.�N����N\�0O�������qBOk���n��0�5%�:i���djO��OIj/��Ob�[�:a�X2�A/�=�#���>��3�j4��4�Ġx
�{{�_�����A�p��G�7���#M��L���'��q��]$�y�_�3�o�O�Lw=�%<���HCE-���Y��<�Uo�ز+g�� ���i��4iS8n[�y'pd?���Y0䌙�Ȕ���g�?� c���`�Ę��4��x�厡�������F?���ՑMv3�I�cx�zo�� Z*[?�"V�V��)�	<����h��B3XǰH��7Et��(R^^j�Me��}޴ynT�F謜1�#��jo�����%�i�%{�s0��g����,��Z/:Jn�N��*�5�T�ɯh �ȥp��6}�Ѷ�Jq�*T^:�z�dV���3��H�p3\v�!�n,�O�D/�A�S&���D֗ö���:x���!������7,���x��۴�w�OnEs���0p�i�9Zf�[��t񾕵�4���Y:�Vzˑ���b�-g|��E���T� y�/+'�u���9��U�L�s��0g7�&����3����joHd�=��U|��9MigxսԮZ�iJ��T���2��jzW)A�Ӌ�%��=���`!�J Bp���h��&Z���L̀ �I�6�>]{	c��c�ɚyL��"蚔c � b�o�W�OR[Q���
`�n[�)�/N�����ISF��+f���J`���S`�:'�/�A�����^����_B��-��C��kDzj1օ�by�=9��vC&5�6��LG1e��L�/S��;�Xg' ^�or^��;>�] @`���$�-Cl��
��'�_J��s��5�j�ZQ~�Aު�RG���H�"���}��3O�K*�,dM|�oG�jx�9a`��Y��=���9�1V�k���en�tF{7-_�@�ܑ�D��1���Ye�ta��Q��^;�t�~�@R�F�&�K��}�exŎ�d@nB���7����w�>C�J-j����$����5�o�нL�Rck�ֽok����v(�<[thWҼD�w�JK&�h�*���cq�Q5�&�Z���>U�8��2y�`神�V�$�u���Gy�rڿ�Cz�Դ�i�z�&�Ji�j]21mV2Iĸ�6��U��L�,��[!ˠ8��UVs�*vi7��R)���K����MfX�N�8��H&�$f��;Bf8W��T����f���&/:�v������Q��� ue1��ڋaZ!������H�;l1�5���tsL�[���`�r"F=��){�L���Z��gD��\�q�H�
��/L�fA���b>F1p"[ٔ`�����+���r|����O!�w�U\ܞ~�Gn� ��Yj~Ɖ �!�)Ρv�͞�����{S�6��z�p�.	����y����gm�����[(�A�p
��x��5n_�V
��s۞蠞��{v��.6兿�Ȏ��`�GMq;*�4ĶT�Zy-���f��?%[���'���sZ �X�a�Gk�B��2cp�4�b����!�5"�<�r��6?6^�&#�ߙv^(|H�[�
x`�䀹PL$�=�bv�R�i�y�<���P�g��!ږJ$r��EG��+xYSZg�Y5��A?<e���8�`�V��@ߕ�)+��%O�Q̯��	�:� �����0�o�Ӓ����?�lN�O��>��S���5f ��??}��aɘ���⡧�b���Y�b��e
j�ʅ����Y��mp��UT'o��6�W-���+ �_a7��=7l�]6�<+'!��2C+�R7b:r��G��l!n��ۥCo�
yי��j_G)EcTW��(ᘰtD�z\��w�N���+1Sp�A))S��k�r�S<�~u���}z	���(�uX�F�K��[)�,j��/� a֨�YLK1�>&gQ�X�8��i�;z��r8QD�zE|��:ΉO�!�ӬϞ����'���;z��	ٷ`lR�T�)���t���f�ȍ�W ���Q۽*%8��5�4�0�U�,/K
�h-U����w��\��H˩G79�Z�*/�e��˳�v�"@����,���L�Sė)4����j+�=������x,x!�@�5+ɶ���5�x.����/rc<$���ح�U_q��>�d�y�n��!zc�7�O��#��qԤy�,��h5�Vs�L���>h���-�ђM���@�����_�ٮ١(�΀ޭ!"ܕ6�	�ً▷X�BA�Z��?���;���X|�ˎ�����O�cT�Y��T�V�������씕������K1B����R���k��'�b�C�$�$��� E���j7�4�U��W:���8������M����7dd�O��v��H����.�'b=���iYc�R
^zCm��&R�vzECo�GX�� ���s��C�K�ě�j�P
߁:�W�Q����33�\ΰe�ov$ΰe.>��M~*������Zn2@�D�AL|��#��G�/(}Vd�w��޻|B�@{vf<� @u��6��	9(ꗓ���X<�An<�����S}	�B��QFy�ӧ7~� �o��~�	\�j�"�&�k�+yũ���5���T�o��=�%��P��R������Z��/�!�Ϲ�me�uJ��aN�����"�_p.�)��*M��N�[����T��E>5��kX����P���]�~=�۩jYA5I<0]���U�Aa��E��z*P��������iJ�$^���������������&�g�������l�GU˘H}XdyTw+e[Ѐ��ٳ��34vI)E�LB��,�b@^EU�  V�X��tT>�����Cr����FJ�\�19�_�<�1����|���9e�v��8w�C�d0�g��Z���֙j�,�eg��Gb=�����`'J�N��d(~������[>-���.%��>����4B�q���x)j���Yo���G�*�|v[6~���+�JEw����nO>yҸ��i>]�C���k�ٔfdTV�7/J���s��9s.>YUvJ&�)7������J����5aqu_U�zY�/_n���6#N;0�L�-] ��d�K/�����;��5�:��n��+� '���x�N�6}a��b�	S!�ps҃�u�幮C7<iL%�w�+����C��R�� �R�΄�Z�2�v�U�XC�7�;��G^G���cpN6NnJ;p��c4���hs5#[PǢ|�����HL����I�5�:ސ+"��eC���ũ������I&���E�LzʞW�<1�����Cd�7���t(�G�L�D!%E��[՞��g�����<n���ʸ�ئ����^-�E�'�O��X/`F}@Hj>5�c���z=2O�EO�y�!�r��CЗy�Pf��7�D������d�R!����t��Էfi���]�W-���;��̮�дe"����8����P�w�׵���Z�4��y§(녒y�H��
b��#�e`,�L���,�¢K� )]u��9�k��3"7\_�^/>k��}K3�D��-H��X ���wP��2�=0�,=(���x!�[|iLb�|}���NqDv�x��c����
)�%thW1K}�<C*��X�q1W���#c��\������yc���r��P����q�����R!�CE�a�a�����c����O�K�wp9�H�}['�l�:����K�-!w>_�6^�ZS)�6̥i;�'�
�g���M^e�I�ݞ
p�\�D��s�nO�%#�>��LȞ��x�iw�r��#N1r�h^׭9sv�m����RR�q��;��F�mp��Q����q�(�0���\���0��)Vc_�1n��mB)�&�?R�I���?⛱�ߌ��s��æ�=Љ��e���NP8�Dwwql]�E*�P?[�kZ�롃��9�.��L�z4�K(��9\��rt�,7+�jS����lPԽy�MB�փ-e4��~Y�up*0����\궎�v"��W{�?�5�hg�N�<�7���-�(E�
d��)<�����i8R٠4!����A�\�qQ��K<������Q��;�D�c,��~��33�o�Z8�(zZ�Q ؁k]6`{�HG�m ׫4�4J�8BJe���G�SHH�^��6����w[�����-��_�.Z"jJI�7�s���9�v��TJ�M��V�]ّ��=��f�=�ȕT�C�Om+s�K���z�z�n�V����wY���D��56ۚ_��k���a�M?�D��#��z�M����z���+�d^�U�����o��R����3L���Y����&�ܾ�*?�&Q}y�d8�2���s�j/r|=�"�d����Qg�>7@��(R�м*�-�����l >�U5gX�Ph�K16x�V�oD���N�jȖnO7�.C���vm�� ��i�R�̡6��˽�����w<�^e#�����( !���O��kTm�׋�.<�u��`�yܹ	>�\��C����|�
�8#�xYJ��@_�с�F���$*)��6d� �T�����.����i��"8`��.�E���؄ĔӀ-�eq%�֢yEB�Wo����M�K x�G|hLWF"!UP�q����!=G=[�A��HqG�@O�ɛ �ȼ+�emwR"�(�"�Ⱦ~o�?9�O��W��˽�TO�t�2��&f1���k:���Fuܾ3�^!'<�к���1�T@8e��k&��6`���:�25mq���S���y�w�Ȇ���R��}��	�c�uAj�PI��8z�!ݶ���/{`�}c�z���Y����k�G�W�����n��������P����g�*���q3$�s����)d29��f���� �$]"j�ƒR�G�{(O)���r����=��}�Zh�2{J�����r�1���mlauM�����Q��=��s݃�^��9N!!��IL���l�Fh���!��4�QnMW���D4�!�c��W7����5�Kao
�՝�i󞌑<�ɸ�"���^�l�� �)�Q�d�l7��ς!y9l5qA�����H�C{/��/���0i3yd�a��f�lED���_�o��A��rɓBI��b�9{��~_�B��R��HÐ��HC����������6���!uܘ���${���w3ְ�Fk�=�Nߙ�
�C�,�T>Ҩt���2af���bM+��&�Ί�Y����"#�r �I���(�.Η����_�h����;�o��O��Mw��Z߇[@�WЄb�֗�GGH��d�E�x��a�44*"��"��ַ��T��M�{�����k��R0�V�s)�j�S٩&Z9rI�o�!	�t�e��E%_?a���c��S��r���<)%��=�4+R|��3~X7@hztԈoU%��9�8x:W�b���n�)J�`mM>
�)��¸�{������L'�����*����fa����B�-�3!}'�_�=i��͑�����U!+a����o�2 2()��y�g�Z��,젚���2���9������r�|!s�����aID� ��k��}�,��v�/2������`�׳�_e��r��>C��Ig�mEa�Ǫ�f�KM�H(��6�-�n3��e�#��`�}`J�ML,�bY�=?bEy<� �m�O,�e�!�p�F�|�;���V\�4��Dm�S���--(a�BiZ{�2��+�Xvr�v�M+���k�`�E�v��Ko�GB�.��K[� ~v�� ;!U�� .T�K_cy�F�z ��� G����$(�0�CRO�>��������rqvX��Z��g��zY�X�h�YM��~i��y>q���>^�ɉbX�w�U���U=�E�y��CΎ�b�-,��+l���=��lk�Q�3�NQ��/���s�7_䧋�wZٷDUBm�WY�2i�6�o���E�ﵔ;��d� ��S����JJ� 6��72}$CH�PnZ��x���o-D�v��TC}��]CN
��_����m�O��T�SI9G��c	�I�M�@�=�I]�ݵϥ+-(�:��b���}��mٕ舌�����.7D�3��J��K!�\�c0��Lp��#�"K"y�i9��Ơ��#�k�5Kk����@��~$�d�;-o�A��NuI�3�I�b~*gXx���^�E̔v��7� D;�>}k�*�"�"�ر�q1N,�����Zj7?Iq/:u~Uvm��@q�!��m���# ���Ϳ�+�.�P������'D�f{Tܳj`��?�����Uc<�Ӧ���>�o��6��[,�Y*7�[�03���.F��0EW��،ReY��0+ƾH�����j`cz�x ��� �qr	9�����5sٲ>��o��YO9_:V�6��������>9��0J��~w�i�f��3T
��^��xk9� ;�CkS;��t~_���e�\����y0R���/[�n���@.3,����c5Ц���>��0��Ga���4Y%��D֦��:8����b���_��Ա��55v�+��h�w��R&aK�� ��4�b{�̣�3O��"¢%��I�}�ssz�ze�G����)K���GZw���|nP���������O!����9����5�M�E���);n�\Tx�wl�g��>�+�k�@�!�˽mhᦚ ɫ����2;��U�e���<��#��N0�C�N�0�"���:����t���~"�����hϔ�`i]v𱳼��z-�C���ZV��g�1)�k]���b�aw�� e<Wl�7;��`N<J�T7u��&��J����_�mr������"u��^1S����k4�U@��k6g�p4'T���hHe��g4�� �	ҋ��c���R�~�+���Fc��V������e0I;��	����Q����\I���	��N~�a�Z\�dD�ʍ�qJo�_ɲ���x�KD̴�T�7�}a���ܲ���,W�z�jc���J=FU��$�Z��N�
]��u�wq\�/�e��Fs�cS�Q�@�3Ű�"�̊�a���8�ܨ\����B�l#�SG9e��B����G�(+���q�U��XL��Y6��.���z�sr�U�F_QZBZ��{����#_Y�ܾ2:g�S�w�J-������uJ����:��ټGO��>���LP6��7��D�� V�U��b�d�Q���� Ӿ�T	Q!��ϼ�������BS�b�<t�6tU�S�a����86]�v'�gg���bO���������_�0R���,��4(z��c���B�9~��ʏOa)�[��-�3�9�<9�C�beu&4�U�Z䵠�����K��{<��Yב�B�~�[u=�� `�PN��A#���YK�N_.�Z�%S���y��,N�Z�)0����D��Q��rU�c�PB1�ΑX���A;?�S���>S ��=��퓣��e�*D�ol���;B����^9�$�מ Z����������#T0� �!���$K}V�H^E�SY%h����� %uBZ	0�"��h '��!��3 �5Z��9���g.�Xv�ɩmg�(��Z�H�|�:���j������@ZIX,ۗ��0���P��o�Q^����Ӳ>�^J�猅�'�x�m�9ךJ�6��o]bNe!yϔTd�]6�?5��0ut�E�$Ʌ�R�?Uj��`�r��n���l�O�J��2-�4��!Ss��}����4ygI�:�M����;�
�\��j�|��ۛf�zy
8�2�:�-��N%Y�ԓ&C�b�B�����Y��g�9T��U\о�[�����nCA |�'��������K�tK���~D�J�D��8O'eS���?��ʴ�X�p��'�Ґ)أt�+#vZu
� �(vQ5�[fR�>�����?d#��L;D�*�����Hd�--�p��ܤ`0�Y�Fw�ӄ�sB4T�����HH���t+m'.+��N���/�E �t��+��$�3T�N�9�1n���B|��G �D>&���c�_�Nǩ��9]�G#c�Ue[�H��k�t��מ��x�C�0;Qcn��|�%��?��sm�nY�戮�T#'G�t�%��9,���ѽlĂ\!G�6�:��9w����X
>t��I\pT����mN��p@�ւP3�����1ܩ�{�R���*$D���ؼ1��q�Ѷ�y�Z�zd�~SNf^�~�̜�Lr�fs\R�jq�������Μl����A��Ψ/ ׿��4!��z�j��}h��>�������r�:<�]X�U��|��~�p՞��cM·=�i�����G�I�y�w�W�����7�^��^ɗ�����Yn��U��KR���j�b5s�Uh|��q�W�^�5:o�)Z��?آ�HO��]�H-�b�0鷭���H�<:W]pF%�?+��K-ht��rx�FG�ƽQ����<�~��巯�*�g���*	���v8��t/R.�R���0��r���WQF1D�i�aB �^Z,��=�;��襑e��L�U�f#	���kF;�;�g#����c��\T�� �hի)����^R��8OY��vr�	�V_�����f�/�`3�;��=3���ƺ����.��t8x�U�K*��=�M8��zV��5���G>Nyn��!���Y�X�^�P�\�lD�r���"PT%(�c�.=��L'v=�9�0$��<�ؖ��G��t�׊�;�$����2��r�,���p�pS�`�ToQ$��=
iJ��ͳ���M���p�J>�A#����9GF~�����D�<�8������w��i��m��˭gi�Ns��/tL�T�!YX�v6\� ��T�pQp�ƺ�Y���=I�:}q��z�b�c��=fl�{Y?���f:� ������A:���U0�T䭚�l#zG2*��ǳ�90c�۟Yfh!�k&�[�K�T�-�����h��;�#~l()�$�}����wf��M��WP5K��NC�5�'�x!�Ns�c��o�_��N�c����J}3 "ư-��7YQ4^Q�J&a����S0ђa��n-{xM�(�ӭ�oE��"�è���!�~:Q�m��%/�7��~��w,nZ���e��]'v�s���(��4	���?dG<�I����׈��TP��r�2)e[�e�#���')f�Cu�8t��`�{ܛ�'�3�'��j�0�A����s��:E����fڊ��/���e�܃�9��\��\!wl:�h���b�u^���z����&�5 [�m�J�x��_�����&�*�7��c�U ҪI1#�)�>��aVq��,���Y��409��)zo�)֓����=�a�QWu�cp�����+.�o,>b��'�ѕM�_������J��4_�K�*^�a��;�D�}̽A�V�~B�x�	m�x{sV�F�/�\���1���l�<��i���X�DO��Rỳ^\r(z(l���5��ӧ��q��$��G��79�(@-�;;��/�g��_P<��W���:Q��@ťI+�RIa�u�f�R��
h�+��Ѳ{=AV·Oy�����l��(��n�Ý���ٷ��xn��uT@����M6����+~�P�[H���m��- )@�D/��Y������UezCə�.r��.�6��%=6�g�1����F���Bϙ�O�iM;����	�nq������S�D��뀌��ϝ�s3rOt	�7��oZ��-�Я���@5]b��13IK�3VO���P��4r�p�.@� ��`as�'"����]I�BӚ[�?�{.�X-�R_ԧ����g�-��a�C�L%�+���%��Y�� �+��O�����{�ٵ78 �K���B8S 1��ʅ�Σ1L�c�P�7};�����ڂ��c�a���9�ׅ�E,Kz��>9�#Qim��i(b �?�4Mͭ�'�����+e������J'�C�Gr�+�X����U��5�wYU�ܢG��h7Ws	8O�����a��&��ae��2��Q2y����ם���e�*DO���t���v����E�>��d���(�xy(��\5���<�(���#(�&V�ݑ�d�}�s��5/D5����=���c��C������
������g��xeX�t�^FS�wP�7I8e��E������	HIU'����>�u��Ey\X��5�p��'^�[9p����� �[������4�e�����#���t@�a��u����lp/otڒ�bV�^���f��6>��#Q^k|ȯs��L=���/lV��B��?����b�8+��_��tZ��[�V]zr�A��w7��.c����O��w�4!��Uc�K �ָx���vmq������@܇��;����V=�Ӣd����B���ˢ0��+/�AkA�'�zٮ��2��"6č@3Q�=�����62����\�#�WȅZ�J��+���+~��U!��������j�4{����^�f�����W�K�䨻���2���YI�n�=���љ��[���{7�T�,�mt��g�*�	�I�kf�����\pu�;���4�
��Qr��I�o㗁��7��C���� ��U�D�2�6fux|yڬЩ��Zz�D�,��\��n��N���5P:n4��i\�R9��T��4u};��cզC�;�GC���\�˸�RZxX��[�9?s�̲�84)4�{G�C�W4m	�4�z"���C�������o�õ��b�Q�a�L���hz�5GP�}I2]]�wO���v��3P��t���e'�k��N�8��j5�Ÿr�%���mW5���b����tX��2�O0��Х�TJ�z��sm*�;E5��T�
A�����<��ʾS�}��`Z�����bȧu� �?� F/�	����Q�c��v=�.�«ͪ���3 �A�ƹU'���,����C|Te�>G���ǔEyD�N@<}��{ Y�X�c�غyu�D�W�N%��������v&���9��iD�a"-AS�*�B��6	�=N��Ujt����&9��:��!��ԔDS��V��A{r��Uh\�ͼ�\+�A7?�;=߸��<$f��eF�����w=wU��~��?J�.�q�}�PH�;*�(����x����u�ևYN��`��"��G���I�uF�ע���e�EC!"�V�Y�E�%�eW�H�>�����T����j�t�cYN�Y_~(���P�ݦ;(�z��b�v�sՄ��tZ|\�Ϡ[�S^�u�58���`�u�*�/��9���%�@љ��$n�"U����Nn��0f`D�W���Oj�8>0�%E|�$щg£��J`���F:Bg��K3I���g��j��==�6�@_�5�A��u�b�p��J-E�E�J��"��P_1�R�c��Ͽ�ɱJ(iJ�Ulxx��6{���;b����H$�ť���;�9��k�$�p�[j��=)vL,Y���32	�����sҚF�ݍ04%�L�QϦ�N|��F���Td~S!,�f�U��}���[H��y�X���8��ѝ��H۶�<�ӯ�2H�t��"�qPR�~���a.7&�ֳ�X�?��]*:�_rK��h7��2�0���W�`�Q�,ᬢ�p�o�����qP�9L8�Ϟ�5@�J^�g�?n�� ]0��3�O�m�p�E��l'~}��]6'h�ss���WF<,���r6K���q��!w��=1y��K|�>N.
������L׵����kg�4����ݘ�t	��_36xI4Yp^}tT{�-��￈��C���Q�|�#���1��覕���daw ?�q��8p=@�'	-�����w��3щ�4'��݆X�z�_��� �4nU��
��;BnIb����ט�Ӕ��8م��^ % -�F�P�c� ��g[YyE�[�,=a��\l�Q��vF��}�w�9�u�(�X��9k�����g6A�_I+)��ݾ-�\�aM�>.�����Dl|��ʻ~�'�� ��j��-7d+R�/@w�:;��L23DS��`���}u��[���K���.����)U���/��ȑ�O�F;Rw�6� ^�A��9�2�%��g��RN����#�/�}`�h�a�	�ڧ�1l�;�V�| �U���ؾb�;BL����U�&/��Am[/����,o��c�;��u����se����v嗽�H�</��y�0[I�S�r��һƯs�.�i��V!�9z�>� %`�UsP�wc��_,^K��Z���R������"R[�H�B:��~��5���f��C|�����s]�����-�a"maF	���,PL}�u�'J��p����of�׎�����tM��/	̛8s����p��h�` S鵂�/�Z�W���;�ر�N�!�U��&���Z�^2�P�󽡷b����s����?����	�/ s_��b���zT�{�H���M�n^�
���*M�16�ɏ����+��X�9��jK5'�I{k�1>,��A�2����t�*��vv��̓	��	��CSAYפ���m�$�����Zu#�f̱�����7fc���(]4�~�٫K#��^i޸#6�`Y����nڠj����7f����"Ժ޽�����&�E�Ϩ�r�=Z�>��
�ӌjz�^1F�W�x 6۬]�����>�vhz�h��=C{�8�FW�:�zI��*h����yi���1�8H�Y�F�$c��<��/��n`2"���R>�*���e�\���b���� ۲�� �]m��^j���D�U0��p�|o�c��1!oZEO�V�?����4�eg7y����X�˖�K#k�P� X�
܀cR���I���Ώ�����ట�Yړ>�E���@�(��E��)Ѡ�)`��C4�d�L�oq����L��:X"|��N�b�vL�w ����SPs��{a'�=�-$
�
)w�l{g�b^�����R)2"l[���9�$~ނ�r�'fsV�F��E 8�՘�0ߪC�^��Ga�Dm9�"�����j�~�je+Z��K�_��0�n���V��x%�%+q��ؓeh��rj+N�ʒ3� ��7���\�N�Z�Y�N��%�������B6�z��kʬB��y�Mj,g�{�5/��J)A��և`
q�VVG+4����($#�����|�OV�Z[���A�/2��4�9�%��Ύ�W���ĵOj�~)<Jѵ�G�>Azi�2EgH�U)�Kvl�bc;9�^�μ��.�R�;��g-���F���L�f��K������y7s��0W[���vΈ�E��;���''���Ҭ�� C<�7��0�h��c���� ���/�BG��Fa�+�.jQ�_deI
i[��o�u䮣j�[b��EBve�./u>P�oB���@F��E����H�pE��\���
�/-�P�tj�R���r&:"�/�~�/�y^�~D oq�b�.mju�pO�__8�Ɖ;>-�@�*Q"��@�7�A���^O���J����t�Z"W����]1�{qX�ty����4���Dz^��)�x����rm?���!,$q{��=Hi��Ӌˈ���so�$0o�"v��$�3Ԝ��M�g�	�*��@��ڰ!���F&�_���Vu�]�)s��W�O�2,�N��v�Il�8��7���U��n�X���}�:W��d�H::Wv�1;���o�5�!�
�3����.���<1�=��π���~�hp9foen�n����Pކ
M�Q��dMqw������$�t�e�M�X���n~mb2�:�Z_�j́b���L4��9�S粎�3s��J��[�EZ�jR���&��>�B嫿�?�$L�y�X��{�K:��^Z|��\�W,oف�U�x�X���?r��ZS@�<�0��3�!|k��F������E*�L��,��ֽ���u��	ڊ`���;����mB,/�+��0Ɔ�i(�P|Ӆe����Kq�0��F@Z��D�6-mXk�@���������N�E��O�~�z(�:�������o|��֘:UK��D�ׇ��1]������^0����cׯ�9���	ӛK��#���M������;�{Kq�R�>0�Ar�&j�����>,S����?�D��P��:*#4�Z���)�|�.m�P���̄S>�M��~C�D;�
���T�E�=$(�sn�����&��:5bn��={��f�W�N��'��"3�EgDAc>�F��%�aT��� 4y��j��Gm��A�C)��	m�YW�������@s�r)��&��C�A�e��fV�l7M���Ĝ��=�夸qY>�~��Ղw��2����Zs���ߌ�ݜ��8�]W��<�i��_��=����8zW���3����w٭�����q�HAȆ�}nT�����]�<�2..JB:'P��8��/�m�x�VB�"� �1�h˙��o�|�w�F��ڍ��:�oH{oC�d�j� ���B����|�Q�NƒT���_`�$�����,��x�l�4�_AX��l����H;ê�y�Ĥ	V���nqE.;gg[$��yz��Y�Z;�wC��#��}��r���n�����-K��e����d�{�vcB�t*"[E��L\�b��B[tMB��m�U�K�kR)�-f���x�q��ʦk8cN��i;&s	IUO'�,Z�����O4� �@0f��1Ң��o�'I��.TY��4Q�R2{zXT]��Y��>�Pww8Im7LMzHH��