-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lBini1KhmlpoUTMaMNgjqc8PvppDVgXxpKEeI1PAUX+b2nZb3UWhTc5M3h/Cx5mVe0GlF/Co9gtj
E0OwxtGpyuOwRDN86M1wtRbCmqg8sAGj8mjQjlTxORed4RdvWFoDGiMdDGX8cGe7TV4BDq+80vDN
5KRW8ntOxF9zKeSDITuihpthlh5dJsly5uYw45WIARrMVj/vEuoJcZ8P5v7Sx9wWo8ZTAS/vfaFx
0+UCJFUVi0uiiLzgoPCZC8/CbNHJxGHZlQSRjr4FYv7gbqZFCUmUD77+u6E0lQx2XgorpXkClb+9
uNqEkQxLujLgFIosR5+c8q9zHGgSHsGUU5pYXQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7808)
`protect data_block
hiPKv9gJ91/IibVihtraEvmgAJbqtiZRe33NJZQjBKI0M3C+4maJXUPpiEmOdlDkiRN12XoWXFUa
kHP5/nKXJiJj9y8qB7l1W2t4vpirL/VDTRF1d27yc6Nq46m16+Q37GM0gS+5iD4V80FgoPwuOAsw
OcRZ3IYN3mujRSsYKaNqdyytWevSw6xE6u4imOno/SrLRxMEoNg8s83R3el6uuwENmVcbn58OxZg
/bRzTlLgbZZeQx4utWYsOZPEPXXJG/dy41G0NKFeVS/qiVuuJ0LjUazuCJE/q3lTMg5R9FIIqxGS
LQWuG3p9wIDEN0ijF3LsTkY02v3g5eSaWqBnbnvW9O+SNyFdbdOaXVeqYe3vY2Gyrghg4G0TRIwI
ZtX8DXCYUgR0f31P7mxCTytZOklgzqYMime9BLPm2AUORDi/AJXyTOJUjqOra3NR8rID2IQ2Ayli
eGglE3tg1NkTRiWHYLJUeXozCxqM9n30jTRNDqZrEA4h3ae0Afh/KOcbGIbv88ZqNL74T18MNjWW
NLxOSf9yszURJR5K032S+3EfRqoYgf/+miXb7icARm2QKFo5sBJ9zi2pS8eTSfR/5K03CGZq7Aas
ou51R9XmusOmnvL+kMPPDitqpYmGIH7jUJWeJgveDo+Kx8ztOhcHmvabOWnbBSS0HdtRk9fW9Ycy
f+gtNkrUyqxkPC7KJQFYpwzDBJOFr7yQFvymabsU5KJNXAVXrMwf8UCjiqMcFjpM9kpYtQG3ams/
ahC93A6RRBoMXZWgWWt1fL2iRVSsavvHcGmvR/IblsIBhZaX5VhBdZ+Wmli1nNx6ocFfpPTO13Ol
knq19GbpKeYmDCfn1Kr4mECjliBbXsGtUChGD6vJuCO1WacOT693eae3H6kzEuzFweHp0LxmkILv
p28mpfdGRFFXUs0NnwtBrRE1hyBAZuxtLkV1his0c0jDs/stJXENyTLLGYMjfZskIcug7XZfw8/Y
0aCVTC3KFQu8uds7Hsql6TDteejPVmBxF+p2TTLLu81hpQwmg8wzhHxCT51S9K1oQlHdEkRfkZ5m
EHpgtZSEjPvDJr4PtPXfJbSqolV3CPjWO2GvViod9IkGi8K87VG19+MWVE74N2nFQ4s4f6QxTF14
J7fEMKrNHlAUsxzRIpoGCqtbVzOs5z2Taxddls9vQL3P95U+I7IoB6+XoOw9AwoMR8DX3wpXgig5
9i2HoOZxtsx2V8HpFo6mngkXCax6H/hFnm+PzAKXy88RoEv9Fdir1Uy8Km6/+7o/0jEJxGOvBkLP
8x+h2Hr4TYV3mi6/WuqLeaxx0I52jJTik7jBdcEFZksNb2eih0Ihgqc5yW2dep4rvbFWv25Mol5b
1c0NhPwxLOTQdlyVW8QBl3cbDzlVJsQKcnZqXl79nmmpoAgI2lPlYmoM7SfeCpkt+GxNFhUGgM4J
mbxpU93y076PCYJYcb0eKEMKpFAlKichwjCd4+kwm8GHnDB6iZUgv7gglEfMl6clfb9B/xD//tud
uCIre7vMmw3W8ZCGQKIqO/Scjx6g0XMvdR/sa01WA5UvNh7Eyf8YfuhPoMaFOGFkWF2p17nLELcU
JX4AHKAEhm5S1SUTXVS2W/V331f/i3dJbuzM/FNtdgOXMecME3/sdnZWuPotu0k1mBlf0sphXSCV
+NuAad6LQwOFTIRE4aE/aHkZqAqCHLDJnvt+w7Kttexo+Q7nv1xwSoNCKrKNhUbqL2fNkb1p90F7
OVl8QIsq1ArcnRxMYtwKaNfLfEBV1xfquAjlOZSn5/oYjy0RbfhK28wzA1cuaORysZ6UyUNJoo3Y
u2tTIO44ywnTsL1WzYhEVd+7Mg2m1sYxxWYJ8Gydnm+a0+4aF12jyhtkrFGiEK3Hs5c3XbyEYzZR
KpC9tsk7/X3iH1uBRiHVXdANH8X8DFcT5+wr/cZayQC132ih3YI+iHad1mCK/ItQUoUrsawJB8Di
MOobW3qCa8LIsRjLaRdQcDP8J6IhVSFOVJj+w1BkNt1wrBUnIcUCzlRhxX9zjx2DNH1u6eNo04Bj
o9stwJHxcanwx1BxqjzYshyFDiCMHHLFCvrql5eAFaRmD79BclCmMYcu9MjfnuQk9MWFHmBA3V3x
3NFDgnqBYtsrgccd8hgzIYlY+yBwDzTZ1Foi9M1mgHMmUivqC2oVmQzqDrXZW60at5IdNkbPyKRY
kem6xWpiLEj0qo+KFF3buAuh4dwNH9w3ZcgYsGuMgiHe4b4GQh+avhnkFvP+1Hac1wojGy1TS8GU
nTWDyNZLxsUaMNQeMIWp227gyauNePEdB2mMuWgEU0pxgtQDqKazs1OYeWSr+qw3nvVJPv8m/HNm
Q/RfgOSxBiY3cP3HQdQQn00t0AEae3JJPWSRNpp5Kk2JckF5jioSUUJUiq18sZxn32Ml9XDtCvsg
nUMxUdByloQMXHrdcnLfb4AofVy1JxFaY+HLHORKRj6akwfVmyGSi0HWTqswUfcosrMuFCQcDbNh
ufk1p5rhlLmVCt3bhkPQKYX65308wgQyvFdKAurAs15u0PnqaBAZDfRVeBEEd3dYXpmSMloYsmZd
4fiKmwFKEPPnfY2rbIS/rm3oKMpCxz4mQkZhvv6mIw6BOUSCW0aNZXGxIwhySbF7NyAlBG5OnTBg
Es4nct6dI43ZMZiiosayglPYY4ny/2W7xYPYw1h4UHYHHeaKRv93A8QUDp0SZeUJOJVVHnCQA0bs
Fkn4xYWAhSNzULda1BUKYbauoRG/z1K2A8P1TRV5GWKE3DBsW3rfT5caycmXUowWblxtpWVR4g0v
4sD3utHb6ZwnubKLelN9CIZH+zdsYuILKSS5BT2yCce7rqRsDn72uTdstOiNsthc7+nj3z+H0wfV
+91bF3ZGl/Aw1dcyje55iI05QsthDkhjRd8rFt9vvYSDcMjf8sIBdmgO4oTiUhvuyyajBN1IegKA
MRKKA16zkHlUIvqkD3cvv39bXvwlO5OmC6UVLgQainSm3FzuqTukp9xvPXYNA4Azicfh/gZbFy23
3zYva6QhZTe2FiicMP2iTAn3/EK35J5ZAB0zHvJJc+Djv5NjGIvady2oHUjBLaROPQZ59CCIYMYl
0sKtcIXzLsl0/Kg7caWdJRwrUNnp3YKPk8MrI4SRtu78kX/G/mGXv/pnthSi6VZeJ4DUbdeV+xZA
KzQnfgKMrONQkwygIe+FgIHmHlx8AucimNsJaZIEz1L6XTY2+77ctpI6dal2YB9JcqpqWgnmRPt5
FLfdwQ8PobT1CIYcH5wr8EMiOZTUzfQqyZT0YDGtfm4TDZg/geSPmVKqeExsyjNcKUnsiUb/T8TE
/Ftp2qg8Pk3iA1sHSF1rDHun5tpiE09IDoQjQQaSARbZxl6yHhKIV8TjDvGx2BMtXDc/8tOezKdD
vkJO6+qiDKechhKWNUrzU7+tyCgZ695rh7CcK3jm/GjDg5p5e7iz2n5ZohszYFNpZKSu9Sf46NIE
of4kSL3Ox6H5jD9HcBqU4bJuhBW90RyJwydCw5dbLtdGW8TO5yHERYSAcQY7h8eeiOGxU5sNetyO
k7gBqDBD/ad5LRmu3krUFsGUa8uIqlitGiRDKoHaUwYz+LeyHCQm3Uopv2TT1NNwstWvYEiI/LXd
zEVFpAIiz1AEmo4EA54uDNVr0Y2OAMtHS1nPUDHp4cl7OJcYwlOjlDrjnSf7F0z15IH68bu0aowp
ynuEF2QSkvHRNHA+2W6Qm+ezUfYgQpjZ/Xv7L+amP0uLT/JpIWlkfVFq41fTOc5LqsmDDJmR9K/d
4wKQ98klbC+LdHarDPdkH2Iqd6yZbYKbqrYrQaeQeiSP3V/L6B9u2LNY/aLtIVruoLm0r2cPz0ST
PJ0KPaW9LXUrxU+sqH5itW3uQJSdbF+WJAXfE9W3hi59skrPbUXgOBJqdu4GcdwCCNLZJx2IOI4C
3QAdokxCrbVC6XHiKXMzK845t4948GCJ8KCfAaEyfxDqyrl+Or1e7KUiH5uC2IdWmT5tVEatbN0E
wR+JobIZLABG4Pqex9snBTWji6QFM4mdh8HGpWfP7+g7Zv7MHDRM2rhbMuJNd2nYqjknsLnH47RQ
DdzrlplqifljDxFP4ckviab1JL2wLcJHkFlZbQPajMZXx2SQtVD5dfLK8c4tGJMpwl7tAgrGfG64
JjufgMrYkA0DZXoEJVrz4p7D33b0iz3MxOWkQGVHTCXcUPEtzMl2qC/FgXJsKc6cL2tv57VK59p3
7o0zP8IhHybn4tms72VbWMnxqQztrSfrMSkVNkvFBimhniqAKh0v32w6yIbzFF1f4e8JjgdJ62KV
rGIeivkpFAGoRJnP460uzkTqwwW5xCDGNDFAjlKpw3FUg3LxJ2vwGr1H+B0JclmeUm9H/ZESgoNj
O7mVFUbA8Hh+/Y2QjsO059jvYPqCyRYvUVCIJBDQunn9Aq3Myb68pn7Z9DxLLZ+ShkjpluyPXcin
aTuSBsQbrDcMFfJ+d5kv1ExyAXnL0uCzw2ysspV1YbEQUIStQyiBFOfyobh4XOAnGjN1UAJL958x
WHyy3WB2z4WGyC9YOxOgJ+GbsUTRR7EpeemlcF5JEc9oa6XXDO07gi4ha/PnUcXye3uxSUAuY7g8
2J2n/WppVTKheKNNXf004PR5tx3h/W6ygvVLwuyaKNNSd0vLzvuyf5B9JO0WC6befm+bOA1ySYZV
BfwYek1OMURv4+lwVJDc6c/j4y7VXYG2Qwkb46U2g1Nc3X6TeZtUi6pgEa0hS66UYNRXsUl5Pyqb
T+xjtXmVb09trezciVSImP+QepOIDKIFX4Zc3N5/6v6OkQ4YZon3+mxqlKMD4arHxjU1X/MN3R7L
a6AOWKwELNxF5EmWJ3Bf2K150NGaWtEGSfkupky61DLG4IElmLWYbDQU2rgniYBgYwh/XgHXBNvN
vILKcawRIuDqktsA7c/hhogP+AEZ1nzUdl3jxtuwq0Rg/RLw0bVVgS1FTO2rgq1xLCVZLOQoFBBW
ovJKaHRMtpFSbti/YscDKfnq0lpUcDfk0UGjZ7VRbFw5ASmcD8fMhQA6TBLM/StDQrfLSGU8TR3H
6VhcQIMFJzmwQOU9j+x06e1S62bEAL+w53eygTc0FJ/8/WhkA0OOrvB+Faxr0injMhQF44aHKwpl
wmJTXCktZM6Y4ZqKUPbIdO9Mkz48RnphfQyyCYeyzaIQN/Q91TvuZGbGJZUH8HaCG+F857Z8jEVQ
6AephNg+MrolZPxZIE1L2VJDnzutX/7219qQZXt6VR8/fb2YPMoxjSfb159HwwUAeEuPpHFPDn3n
8omnvtABkqrq8GZ3SwfFf0M8JFWGkyv76zr+bjLIPZShUSAXVn14Do4P9JP/VGnHSudk+LHA5R90
oq7B1p3F42vMrAnNcbVFZZe5Mz/hkfS9vHDg+0hS3mD9Ably/sx1XQjcoN8xbeOl3B9VJ5UuEiWu
kRZMq/UoXf4KEzLon6ewErfeMI1dF4/EcqCu345xDb5LVEDdmoxLsIQ9gcqxqfcxEqIJmsXiDzkk
IchFUveAgcmWGzjhDiDE8QR9xBFwn1Zs0NlkPh2+SDZQhkovqfXfF77Wbw0isuVIWp20+a9Vgsws
GZNooxBWX6OgTx4LD01cBpmjvm5P1R368Q6DUKLGPn6AbwezZ2Bde/liIeWAoZi1rikdXCf42g7M
WVzhYhpJYVhRK78gGUAG639T+6lS4gr/IaAo0X/I41RR+XJWBw2uOlJvIraXHulCG7am9OzwOmSF
fZIAjfOCU945sTiMfsCgboJmdubdBdFAgI8jODIj+mdhYo2ZMG4PykEn0qKk3kjpXJ5BRAgw5Csb
KA1JnKLdYHQtU+HVZIzzr8zgML+kyaYXcv5n/47wDkP+8eh4CONDjY0inRe6raJbGZ7WvJzrYa4b
4pcR32vdnm1E86k91w8MBKkyCjyc3ndfEz9Nec97pxms8U1o7Bo1gGAySgLdqOhbl+srcpxnSRpf
9TsFC9RGIlObI0X79v1rmp8UJWIroZlJg52MQoOiHEKUeDUqK2VQNQLxxBzTGhs1bx0063Mi6wSR
rCG69Kpor5HuI4Iq7byNCPZQC1CdX8ELbt+uetow3eAlK7Mtq4Q1Y44uNqowAbY9itg5XnRnpOxi
gXOBVwc1CSOpGg/uScf+FP+pm8vwJOkFTdq5KnOD3vELbeDQQx+fu6lGDCPk+DTqkR5Wam9EkvFD
U6cFD58Z4aNTXflwImeEo/jcv4qXzLHTHjRMNR+zWgQo1ahRXwC2eXvuDY9PuWt7rD8NQOmhXzsj
R9/MnyXlqZhnmFp8JErxi/AgAYuuD5QunPS2mfwhnxZ1bkeycnQYUhW4EYfRULoBON9E03ZpfmKX
ZaWLTtE5vTAcZmDGyO2LAh0q201GE3oUZEzlAQXfXD+CXvHgAW1oQ6a3g68g64nTI2bK2WMGCwd6
AQrrUJrP4YOXpdnpwhylFPXFoE61jeJ1h7zpnlPfWDwedAiMLW7EZYIllHmOrdyeHxO3pLpoPhvX
tRM3tOfuuo61fjU28PEXeP0AoBPDUGjqdGxeNpq4jnrVg777rx+iPCJQ+3Kil4nIGsYZTAlvclT8
iQRJ4jnTKA9PMf4GNB242qddsCgfwygNN2KCq3ZGyD1fYP2GcRyuMTB9fykuowWXoWot+nOQ0MTk
KSXm0ReNxATrq571/YETYR5lYJ6WOBJB1Hwn5zYyEODWO2/R5Y4c+GSQgF5IMrmmCw7JgUmW0UJh
yuycy+DhXcA76kErYLpup2G382ENEMsvJXEucbXiW3mZegRx/3P3Wc4tSfv6zBabTGvw8E2whihx
gHlXdEX5QsdIx8yKnblEN0ly2AG7Qmx53YTrxotTgzHB0WLdd3zl8RdiAaqTLIJiK/XYnsuhpKfG
QighGVGjUhZoSIbJcqoXdu+1NL0wBnBmyOzLBzxDaDvqiAmPhNsGToUxCNp+zkyvcTPBZNxeFvxG
FcfUGLXOv8rzctAJfa+0HzJUODmczqSpsvzIRaGxJKXBOrBrzfq8B/NbJO63PKvifQtDqTuJwUws
9LYBd4yhgzvTaDUnEyIldGpP8YfAdTVHsNi3X2t7U5AzYgoY2G0StDi0zrCa7KMiP8m3+fL8msj3
itoKPIr3pQ9z2BeXdBnyGIDEY3NO+RrGBrk5cCMMhLYPEagoq9GevjHcnEYZWGDwzPR6l+iXZKoX
axpUuI6T+8PSvcg8ICjemejhSF1tnIGwk83JsVLcq06WYJiwFabyjUc+hyD22KgzXFL2dWgv0zJe
NxUF/SEFIcayfxkuIQqtzn7ejc7mLiufqfIKodnhdrWGsRCHocbrWT4hxK/IFLPTDq6ztbzs8g3Y
YoqjzQlE533lT1kHfDSLz3c9lNyGyKS7LYRsnageIxRh692dYD/Kh4cG7g/h0ulaLyTtkWwH9jA7
g7TnUZt8Zc4DTyOMyL5+3Uf1pegAZ9MhqSsD+UR7slgV1OdXZQVc06ft08XKNPvU0tRqqzD6A9Eg
b7gCqrwcrR/gF16jooK7NG/4Su1mYSLyT/fVr8qNXsrJ7s6MVuOBRJFkHSOJWY55Y/O0R7trA4pZ
IJSKAUGke+hidFOmHg7lARcHxmDpehYGJ/i6yPRRjONo6o5UQEnfdWJkyjNPYWDGA4fV1sHnMfjD
7JAfG/3F+5s4QOCYTRPBVQwERGi20+ovtPHEY9FiEvgel7U5g2CIS/bVTyhyBM4MbWSyjo0LOIWU
coJbOQn8FwYK4GdVvAoZXPvR39689fDaRqKHih2TmOWNmXiJHomfCHFCj3uqGY6rvbVFeGK3Znk4
pHfPVpdoMmhBmffrGnE0tiHEO+P4m6lNs9NWOeoQ6G2XWj/XVKKJelNF81T1oH5P3jc5DZQ+oScu
HMKu1tPWBiucMXX6NihWob4DV1gNviichvAQ2JJy44FQBmOAPFmkM287oa7lCcrDotGT0Y2GJMRl
xtuoMEZkHJYlaEVHQ0nbZn8oGjcV8quGvqNno5FX6delVsFCzR1iDX9AQI3GIHr5nDXmcP+4SBBb
KXrgR22GsdBKAgpKj9HfmqJyePxDHW+U0qh32XGrD5f9y9KZoHVJ7e08qES2E/+5h8ZXtqfNL8zy
QRVBTvxFs4pQQ7EgGBi9pktpOQbFJdPPKpVo9O4I8+uQ+J4pr+AFLU8PZ0NxVjk+WHbyqffOLsCZ
fa3NewDpyLnUpDALtfoQ9M1xhXNsmtVwsqNOzeSQrz8AYS7INQvxrDbWj+qr6EQWxdWtBCl3nL0R
vd8f0vhnWqhuRBqkP6SfG59i+b4/RWkLjvkOQI+OGNJ7f499fPgRtvwFqVIY5TUcQI2tlvI/jV+D
YiSxagS20R9G9UHi5qoefoxjQJVTyPYLAp4A9c54veoVS5ezSohE2/HzFxOkSPWROgb1luW5ZQVM
USYarNSMoz/b1jF/7EKMimZwdgjxLIiv7LDr5pIQtrtRGEla+Xp856qtnx29AKY2Zzq6kwB0TmYW
atO42S0l5yX1ZCb+kjb+U4IeCmg4tTq70tMHT7cwxdMdcvJaZW5u9jvkHM9+C8ylvdy5Lriu917V
q5XAT2yG8vyx73f94GAQd82IxunprQKNQXa8BPO2oQoQq87xCEPJJZQj7ppKqr4wX5Mv9pg0fbi9
fNTgTPYUPh9Pqci2LqYXZNTEKGxJwYSYHDWhaJc14WQLNFoFGTQAq65nmqd5nubpf/RYLPVlPMnt
+UtCQDIkgQEUfc2B47kVy966NZrLemuZ8xvZQ2PmJAYzb38+QhvmgE6JPUPCvsAXHzVSXy8IMOjw
sSPHl9DPYi443VV4SnHz6Pv5yphMr/hnAVVKh2lkdU0Eqg/AZ1iUohvUEbdzk4/28pk2Zhw+8+Bn
qAVdPSoG1z84ZZm1pSQOC15gjUUFKxPCuB9ObOwdOc6vyjaqRw2zNlPGtFHkh85LQBVC4imzTRYG
0L5T5TteWv5gO5O3XfmZCEARoxAjhlyV2Cb/evgL/nf0RAP4IvDs3IW8I8xbIVB7JzAjOQixQeNV
Ev7L2KTwLwXQ8lE/GsAqnLxuORv5BRyoxdx/L5pW29AsCSupLzxlePqfj9E0j+3/tY0zEvfhIlG8
5U/qklnF01IhUpchawnlSOg8gAV38mBTiB0mU8FHba3f5YvLHf58lHU6tjyGB+cavedPsnGOQg4/
IZmXP0sI6fmwhXZgRuTym8XEP5e2x3k9+Z2Zu0WnXXdLd/UoTbNJRkV3EY1y3+z8j2u2aLRXphhy
loKQAnT24ro3pz4c7qac3rg8vieXLLKqHDe5a96RgCGLQ51ajMIT75F1ShjIQmgTx0wlyWbnf9PD
eJztJ3/oqXI6qrjPylDYy/kR1DiACSAFgCeM/iVVF8730QX2cXubtzOfjjFhyd8ABqew8nXfCmQe
ATIVPxhH7j8L/au1h5OhD8EgQHxXEDA0AqDdNvlNlDW7CEO5K4YKLpREQy0Qq/3hiLxjWeije8xF
lk4ToAuR04SZ2zeMOww7E3y4oL81zf34flhsE/m4ASr0V4T7rNyEPj/u+NaAN/IHXvh43dZJ3xwP
JWAijuY0fMhcwV8mhtgPxG52XMpVbkfqatq+fDN+FaYInJJDE6EYYitVLXTSD8uCIwzOYrzQbaMG
w1cLx9dN/OUEDfeMEggOePXerfHcAO+YCUweUapylySXeu5XGsXODZg+g7QjecNyaFBBP2WjwhCd
3IQVdCFr0sSlu+hnQDy/b89JZ5r5infOnSO8aIV18K9aDwfG+LB6M2wJghEczAWuTerehBjohAT9
8VsEcjMHZmBiMY+3vdfLdC7Y0waajmtTY9VzvfTIN0g+FPrhMlvLyNNq9puqd4ICK3yxM4jhBTPO
Kv2BYqx/gG+UwdsBe9PzqDqIitHPORTXA3gwGu9qBlUhsQmqjuDLSsEpi7Lpux4NpobrjgR09XwG
J7KrKr7lZKlHBB5REZl3W5/ovL+GPPiGQzdgtfLKtPRhuKUjr5ROrFoJrlUYMg45GOGP/tML3auf
InpXCrrprKvGMbN1wg5NL3BbMh3LIRqs/AZP5rKTlZRp1Tecri6vNBuJfId+Lll+Vdt0N+gI1axq
Y1daakSkLwDi2TAYzLObELE5zIUpyHUcrXnMcctZYWb4cQs+MdHvR9yc3BxaihPDSHHHOxxUl/1B
jl+FneMsUf4Eo9HFfpuEtYwIfpZHFQcrks+jV9nyXvDUcn9gEfCAarFQ6CrlXcj64SRCKaRRrvlc
dOtRoKig4lsq2YDVG9DAFx4u+BwZ4cs6XgfsAT7CuKsWUIL+aU9pqdBl1jmN2rhlr9hdYk/nt3Wo
g1ZoHfdMFkK85sPqU3mu2joF51p+arIlX2e8o+8taV17xC6ORjM3rPwJENZ9uW1pvKmiRcKL6cg=
`protect end_protected
