��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ��E�[2�Fg�{�%�I�,w����d���y~:�E�tʓ������o6S�׋k�(���XDVe�F렟"^��ä椣�\Nic��>��[x���bR��c��P�oT�K!�4xx<yJ�����Gّ�ش�&�n�u���P�I�χZ3�-�Z��_\�Ư0�,�̥�ha`No�s�
�c�d��s�N{�[����却�x���?�pQSG4�N�����������z��nk�M5��u^�s1����^ǒ�~Cc'9�{�Ն�bH٭�����P��^�i��u@��	b�\-������F;�&�Gh�g�;D9^�/紐�co�83�o�a�c=S��z�Z�`�s�PYĈ[�K�ƛ�>B#�x+%c�8h���C�'��?c�uF�|�5�">�b�fY��^w�f )NN�Jݻ�z�-�B�bC���\w6k��&)0�-�����^��]u�8�e=���Xt�q���<�]�d6�a��O�[�㍻%�Bq�]�л��[��d��F���8�ί�M�U҂~��T�W����tY-��y��T��SNd6�jG�-'���"xG�"X�qM��JMȉ: ��Nm��jr]z�NXg�
Gx�AT�_�.�k�����))`���oKӮ�&�'�8�%x_���8��qG���ɺ�޽(�pO+<ķ��O~���@*�҇�7H�0����t�@�^�{�R��@�R[�*���&J*���thh��c��D�&~�����趣�=��A��)��6������Δg���v���G���xo��IE��f��.�#?�����.���ֆ����_�7����~�藳tN���'�l�h�媕9?�$��DF?� ��?bS��/|�n��!�(�XAQ����c��5B:�x8�:Z~�xX��6�B��s�v��:�R��~)��n���U�i��6�)�)>�%�9���n������ͽ7�!y���Ќ�&AG��m�i�Ў���)�W��g-m_�D�l��-��-O��0p�mR@� �^�pZ��ˌ�@#	�:1�Ov���&L׉)��v��|�X����B��h9dKa���S	b�_J�T��*��XIh�Kd�F�=�%G�Vփ�2V�&��ֻ'��пQ�wH�eA;��H�l��jE�$"�t����=�u���~b�~Y�z��Xq�isO�Ĉ\O�V�]ر�L0�2�A3�]]�ϔ E0n۳��Jb�ϝ�׸�x�+�&�X��ǖ����˪������v�ZA�ѫr�[e_�Y�L���Z��Z<�t.�^Gc�������X��.n����gyӛFd�'M}�B �r�p��P��j�zy&�|y$��{�8�"�v�ej��ѯ��=��3G�*�i���"rS�H
@�.�w�q���Z�˚������ΩטG�:��9�1��ѯ߸����9z���[�66�-�U��Yq��6�h�ADz�Z�+O�� �ym��F��A�h�ޔ�G� �
�X�m��c�}bJ�щX��	АTt�\�;�ss�v~�r|���PR3�?#I�9k��Ʀy��1,�C^���W����G�^�fI��7�}�O/�]�~�̏<^�Wg���2�ut'�W���Z�$F���r~�������C\;p{�bC�p@��i����qlhAR��p1���0ԥ<�$@�����~�ڡ�ǂL�&Κ.�/���N�;�@��O��h�W�� ����K�V��3�Ƕ��Jon_�V��|�X��M:$,z�S��4B��XZ�^a3\.�!�_S��W��˘�Q�6�'}����&��?v`:_n�T�"I�z��K7Az���jMI�}�2���kM}�mWܰ=W���ɢU1j2PX�8�D8���*�G�E&I\�U��N?m�f[�j�K�P}�3��x��� �ŚQ`lu�.����	ũ˙��N/��B��d.��y��������զU��זg޲Qu/��G� .������U� �S@��1ܤ~�3{8Pj�( �k׎Fܷ�L��~����@�0�^��=��f��O5O������"v�_P�a#�nM�#�Tu�`QkB������J�Ͷ�����}�z�������*n=MW�ԔAHAy1�:tIU@�-KE��a4"�Ǒ;�?�C5��z�5'oR�J��pcq���o@�R�Yԕ\<YZmKPr�H����J��J��^��2-Y��։�e�,|1e����EXY�����.:�^�^����@F��B0`;�$�f�y>�WZD�,�-J^�?u�����]�SٸT�<b�kV6:�J���Z����j5�_��O~{e�)z���/ӎ8[}/u��Fq,J���ìxn7�$����ju�~�|��y�݊D�����牁"19V͎�y���ݧΤ҄���0��-HLa�`�l�$����#:�X�o!�I�2���v�����f�w-�h.�5��^fk�꛼#��{}L��#�$� �8a�Kۖ&��`~�\p�*��+�❵<����w���k���Z�Q)GC{�)<��O�2��D�lW3�cs����6_+ÖS]7-Oe��f�&��5�$�m�f������F�+�{�I�į v�Uܴ��qv�8Ne5�8�] L2)�1���@Hy�US��P�7ޙME�]�`���;r/���G;Y`mE���{� �Fɐ�BQT�~�c�,�N�0��*3T�l�'?�$^6\G�u��爃��T����<BS�BY�M<�s����'������^ő��X�d {�%<�ʅ�@,�OC[#(1�n^�����L�J���3�y.Ag�F�صT'��J�g�K��ev*��V�<��?������[f{۪%�ϱ5�gJz�Dts���g
����������]��j�Ꝛ�<X��f}!L>��_̟a��S�G��� ��zS/�	�܊�Um\��^Y�qH
��s9<���]t$�Oi�|�2���lf��r��si�<!�-Q��:.�հ0����y�|�m���n��A\s^�c�t6�8��I��'>�-�ϲ3��DFZ��r�i��Έ�r>���"z^\�r|{>�;��<\��d}&�`d���G`�TT�r�qno�+��g΋��-b��8� �.�n��ə�	1g}���A*�\����v	
ۤ�a~�X�~-�`dT��%�F��(�cO-�^�#�p�u��4��gX��P��.3S}[�����Af�>	�P���÷Ͱ
a:�g�m�:^'%�<�|���Gr}�ekMƕ;�T���4i���z7�2Pyف�[X�"�Մٲ�|�P9���th��l�?���/_�����xQB�D���Z?�;�yD�Uĵ��I;֋"���w���w�Ԋ���<%7Y���ۭ�ɦ~䟱q߉���5��N4�aɞ�u�I�<�Ij��,������|�!������`���MW���{[˝g�M�-8���&�s���JEʝڦU��8��RC+���{�&���vIo��^Ӫk ��f0}G�B�z�'���?$�W(c`<'����������y��3�tH�ی��Ke�v�m%ǟ���4!0Y��BO�% �{D�F��f]!���Jk�<�5�1�yIb�b�6*�V��c�HE��C(E���+����\�Ѵt�������\{K�P�m�4�K
�VM�-E�?1&23 '���|�"ӵz�B���f�n��kM(m�@�R����xbl���q�t#54��$mc�X���K�cf={�2�Bve�M���R"�?�4
�v�NZ�,. %�^tVy�udt��lg�;�A�5��F��e�R�7"�C[W��!�I���fL�"[Ğe"Qf�Q���x�L��(Bz��v<��kis�k:[���uBFZ�&�#I��|GH�T[���Z�Kv�ҧ�7�e��[|%h��b�Bcf^��m�����\/.%�`o�ho�`���P���*�h�QY�!
NFh��8Iľ-yOOxe���B(�-Ku�W�ǫ�o/���O��}�F�k��#.ԫr"���&��FTo��@'��@�3��H4��<l<;���R���!�9Ѡ�6�Hq%A�ix6���ε������e���)�%}6�&��D����B��׺�6'zYa�{-(��OOUQA��l봻7,�d���y��fݫ�Q�=͜��mu�QZ�A�3#�u3�G���mm,C�G5T[�5F{�O����vk��;5�+ҧ��k��7b�� Z�au�;�m��7�T&�_�Fx�&˪�m������'��{�q�!����b,^�@({�Q���c'�����Ǐ��qܓ�7��Ӳ��#����n
��i�oԤD�ᕖ@�[A^��(7��P�Ц2�h��qU���B喥D�ce�Ջ��[$�*����w�{ҹlL�`n�[u`�W���5�*kR��w��;��l��	�<$_4��V�� 2�\�>Ƭ7q+A����h8��*�?S�4B�5J��u �D�pF�T�1q��jʣ�x�#���D�Ԥ�"p��=6u%S�/:ɰ�����CDYYB��~��(��?U}�u��<l�J	}z������|F F�odP���t���LC��sO�I����yM���H'x�6ؚDkl�@��N~�?~�TjJ���"�z��⌢뱶J&�[n���j�L��u�=j��<��� +vy�m�� ���Y�m$*H���1ݦ��`?�����dJ]�غJޅ�)���v�֕��չ�廰����Ѝ3�o�&I�$�$%��A�Ձ�I����$��]L���b0�3Z乨�j٨og�i�
�nۤuw������Q����n��Gv���H>�q:�y�}��5��&�a���-[���	��g�ܴށi�n��Xw[�U���͂j.����μt^�%��O!ʜr;�8��AZm>����0�0Y�X��J��W�.VUZ1�_&��xh��L��~�;[Ԅ�-B3.T��c���n���0
���CX7��E����^;2
�;>��&m�"���u숓��	L`�W~_9�P�Y*Ɨ��j�<���#�����ю4��g*�J��^�T�!嵴��諜�=���3�a&X��64�
9y�lH�����z�<�����g�n�t�8�
�hP��� ��V&߬t:"erj�ג"��5S��g���iCNA8	O��:!�M�h�J�E�3���x������i[Q��S&��ŀ�ʄ�7T���m7/�]��ݲD
̳��{�.�k��m𐃲��h�T:K`J�;�� i��d��j� ���m�,�����9`�4[TtI�0���Nj�Pl2	
$����E;{PhM�{~{��T�KX4�+�\D�,3�঻b_>����]FI��~H1��eΖ�1{)u����Q�k�i�O+�m��Coh��M����E��-<��耏��
��e�}����Z,�
J7���\���0C�=ɛR�-����ɜ�����TP����3[�M&�|��<9
�|�+i򟊔rΕ��H�&���!�R|�2W�	��~��|�J�7����X�6��}�bk˾I�>����om:qj�y�Y^��'�]�-#�}�׾���8��r��ʒ��Ko���c+�o#
�||3�����U�������J聒B���������I�t����k��de5��������$�7�;�M%J���䰜W�c����8Y�ߺ���),AU���;���NX�.��%�9Y/��U�m�Z̴f<n��HGCCe�V�90D{5�&?�M��j&=c�J]��"Xd�j���!һ���mK:.���i"�O�m��3i]O�q�0�
�,D(y1�2k��E~��QP�yQ`������Tc|Q7�aT��]�[t0^%�G�����M9A\K՞���h]��lc	2�\����q������5�F��� ��Qr�%�j$��B���FߎA)�ږbX�뿇�y���˙k\-��5o�?ւ��,�J���[��W���{��>��]�?b�v����F?��+�����>$�E�: `x� ����l�5U��У7��;~�]�A�M�����I�b��+4�,k�Z�pI��T�kF���&JV�tp�eL��#uPc.�j���jl�}�9��SU�O��V����_ ۈ��Csj?���ؽ"o���_4K�~�8v%-a��!����� g�OR �"�A�tw����@�l����9�4�
m�g'v��<�D	��=�H�K�j#i�<{���@NZ�r������pQgɜ��֣Y+���U�Q��v��>Z��V�w�TD����+	��Š���pL�C��������>x��~�>6+����S��)*$l��7d9$L�è��d���D�#c
G��ث`N.Z�Щ@�KP�묟�{�┳�yZY��h{�0�9�n�t�_{Z�_�U�=�r�uv�L��o���?*�FiFo�xy޴*�O�s����7���2�:{������'�H?>P:ѮQ�w��[�J�k