-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mhLn7gBnzR9btxWLb70ek5xAkoJ+jmn8sqOunRq7Ys+oReCv8xIamzTTWsfPXNB9gUcqaT6UCZnP
cwdxvqpmekeYeQf1mHfzX+q4Fq1SqKcidNsVYqXHYXmyKrGhg1ARM9PJ/55RIi2oa1uDCPGGWsbd
lE2Bt0X1j34xmZl+45SE/uiLLrr+0eJRL0t8+/i+3AufS4VWZ3H+jNOXHZQB9tyYDBxId11tluH9
JTH0KLAFMKeTssyqRrbdhE9GJ3DBykwYWLPfqdkeln7GSQxX4wYxybNLMhHHwznRwMoUQWIzn4wv
wehoXIVLzVstlgW9hf0voY5CaBQFgmwlQQTcOg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10976)
`protect data_block
YXkpcNRxuGn3cHaAOGpcqFzrr454eZ7Lo095QZrjfdHfsNtGL2wkDt33v4RC2iMtjrnsXZnPHsDv
RWhiLpqdxox4heMIyr5qyDbn7xcdK5dGZ6c3+NI4QDa3adW8h3zgqKD+SoHDV4DiT+fGV1ut7QyD
Te4eR5DSUtKvPAAWbjNuAb0JgaoV9BO8Sxe+A7cUpUeIvvPSjdny9/msmgOxlDz6CCPjPJLhUvJL
D5BOTM65wGVHh91Q12RMAv+yV9QYWc7sZYC4CCQQ3qGIZG+OR3dxwoNwEyosHkgF8VqiHy/XlM84
pF177y/QDGnq8TsxxdezF3OAB+K5k+SlMRv08O5zT8AYL4g6ozalJwmbpAm1znNi9obRaEj3rDuX
2xVQsLVCkZlSxZqcZA7vDYlIvzYjuWgT8FE8jYR8D1hL8JNW1SLUAqNaT+57lbyaChK95Q4g7uWB
+/cfdYKS7BIiswCm4wRmaN4NlK/FX5qWwJCKOu6bs++3Sf6PMyQO//hVUvAbweI2nDWb/k/x/0w4
D7uBCfEE0IsWBo/vyF0sCCiswVoN/LRl/AtH53ZU+71IoCdHBBFnwYiMaUiovhd6xMRSvWqrSH97
/DXYIaIugacFvZgwfMXPkfXT+0U9Eern7JlG0AHbSoouBffg7lwkc7Y/vU27vatFPlhHaBWGdbfF
2A0s+GmrT+kPWDa8lkQp47xEb11maKvAzECZi0iA3+Jml+nkLfYcpnMYafDk8YvHdLfex9NSBNsU
n/1q+cjVoi1oBwREB7t+UlQpMRD5SEhxHN3o3F7j3NV5iawMzzCWPYsQSqzaYkKciwqxSuQXde6y
/FmS0PBKNzSRUh8kAEfRplwgDhg1mR8SwflsLeHfs1cbif5uYNqStuVK34UVFMtWGz6acIMc+IL2
50EC0qeHB0U4mjwgrhBkVeKvO4blEa8S0zqX/AfxfvJPnNHmJPhv8466bfFRtkXVG9N70iiA3JK+
n6myyz12FPUlk9FCG2tzln4NK7vREvx3iGnxNf7M1rmxOeI+x8HN7zbmQI5mdyUWSABrG3HlOloN
ZxPEOd74tFEf6Iob+HHRTdDxyHWWHAmFLx7Zse4ZwbC7iLXtLSszYuFscjAefiedx8VvWheQ02ky
TrludkV4+6HDvLyiEufDtjQnsKnOOC/etp424ZWVdJdZGqmQ3Irhv0xen9XFK99TF7LaB0SCVXHZ
ihrfBLQ9zcHazpKE6h/5PRhKEeMC4e43R/tMS3PcaY8RlqZsiSF4+tUMwAFksZAktOdHKP8vN+d6
+h4PyZNpnPyyWYKc+EsqduJjYcL+rVyE9mjDdCR4aqKRyIWrkpfROx54iJ3LYpTa+xOGUgyqiuCX
2GJnPrFpmvDAaUaHFZsOwvrgUlioI1iaIjgRJNzCwdWhY6c02CTwdktye5j/CQ3/BmHnByPDO8aE
wCF5UxBGGVf0EPdInRPzvZNM0pqiM/Z0gyUqaU4O85MXtvRRnkrZdMZlgXT18KfybPgtoKDZmQV4
hGCuER5TNJVhQqnV1N+ZytVsLNwzbLDCqWg6f5QLCTn8jB6xIfY7CKssI3kSobSbTkLqr/tn8pk9
atNkf+zEIFsTmT+/evF4IZQf7ELd81N6RyuHJAFyy9a/wOVbWQZz/pYu3rV5ZiO0Y9basW/JQgp1
ggcW52yUKSrHvL15nyaA0IjxBRF6TD6byn30dIyoakd+v6p7KDJ0MTvKsWZdn3039owoZelRGNEe
+PjtsSmD0aQtmB6GtzbBUpzUF8OHds8CH3mQsN/I61epbuoES1UzfqhRYzMi9lTBvQwGOralDxbi
C10Lf+FB10nCqf7puEBNRG3n0hmYJqDsyan+H9MkVy04DED73bAMuP3P1G0FknhhgK/LwYBWnyih
s+Q1S8tK98OyCj47bhi4UyOh7zMZZ614TKWBqoxyqncL0ND5NclXbwI1wuicN1OGtnsGQZY9/PTq
mU+KqK/HWGRCy+GvvtVL1uRnlF1WgcY1I2YlZlM96f/vl/td32Rgp9L4LGYsJDeb89W5i6UJ/SKi
W53sNb+e1NZeiaPM8i9IMgLgk92Bz/Q4K/pkeiteWjB1Xn+GKOhYff9zfQeEU1P8ostMdsfquwH3
wM471fDpxfb3xKeoMAAiKXGGZGYUMj80OrCQ0LaPro2So9g6TTdtRngjPVT8YkELLxB8fHYPOyCf
3WSWytjSlMsf+arZ9W6DL/Bfyb55kmxvZJF7Vo/4EuPyhathbRtXi+JHtz30I/jmjKkf2VtGOAEd
k/e2ABTZXXbImwWCnwlf3leT9lIEaF01Y/MsWUJUhaRYBmP9Uftq/bhuuDaNf8GobrTQ5/mznps5
sxUfSBC92q7FDPOO+dkUMFwaQnNpYAsLoByhim2bRDXdqr0g3/Y/a8UUPd+eBK1Utp8yvZr15Hdd
jM38kHvaEIodW6F+ZBW38d/2VqGlMl++mkZFdQRspWZoCrjx/4iOrep3+nxg1NgDUl9bwI5Uctww
gaYOT9k51B9wlucdE7eXspT4XDGNd18kCm3zUG7ggJ0t5WawVyEdZpKo8dHTA04FJ28AKvJ4Zm3I
8xXhPNsm/sqEm9igld5d2l+gwHsu5EnUqKZzNR/fBSIGhJCVbzFrtcckqeyAxcFoJeFBVfpVN9DP
Va88KpKgsDZ1BMgKFEL0haly1gfIF9CO0VGpQOsja6TYwqsl8Wjjazb+XvihO4OkdVRcARYMgu5N
s6dTg2Iug3MRXQoJZ1gbAJfZKZRFUsC9is6TLMmQjXGhFYrssC8Zm8WKECaSg0QQrl1WKBWr3rmW
xqqqPCMTAeeV+/jS8CuMIdhr5xanSJRGgEYRb9KMO0v/coi79GOiB+AUxEwiA4szy+uzmXhOnJKB
44ePZDzNY4iF1OsdiMhBKHhRdCqPC3iq0seRqeYMENDzGMIMdqRSefq5ovbb8AUcRTxQCxYpyO5m
XvIZeSnYneeva7+vNUVSDt5V5mVcL8rL3D/WUsZHTiUrMAGxe3zruMQdj6OIB6+t+M1e4/krouU2
n+FaOI5PTmBqCxzvI+Dp3Bq72Wfb3Vo12BreTtU+SZAwzWhCT1b8bv9n1hOTr3rS/bqK/0n0+CxL
SIWgG4QSlrEY4p1tY3OtX7WtcNVZfOrNLdZy2O7rgBQMrERC3KLqaGPb4hFNXyBF4VH04C2uUgA6
sFtG/Yf0DXda8tZlbIZ2FJl6h436DtaiqGrEf6gkymyRpFWgPiIHm0WKbywbaV4bVU0FQHD08bZE
FlwGEGJ0tGnUNVjH4/JRfvZK8z38Qqi2rSrNGNF4bSCQsMDoobUQysk4IrDilcd4tQJuyGfeJ0sv
SfKV8rwmR1eLOI3JFn3ZcvRmDQ2fFkCEAflJ7c+kP2imUFZAKCy1ymvOSn++SBdh0f7Ua4jOphMB
3I+lP6r+WPuxjEec2E/RCJWfxHhFw4iEEbQNrPgrwVdy2UR0EgWoLIYrQuBpKe7CZ/0FV+jHRoj6
2R4PJYlOSupjv7DjrraDoFnRehuEJGONdi0xyAdGgoytM/aLN9tpjr8+A46IS7jKALmVDFeXv5DZ
zs4XlcC7I0RKEB8Fg5YrIi2jQh2IKSkZJ86GYel4Mg4zGMPpgW0OHYKZlgqxrASc6JK9dvj1i6io
w0Y32mhLScD0BUje+JuooRu4xBxow6B4IPw5SttUspp6VJw2gJCl7ctWPIp9kelNdIHQyY5h16TH
OgKO36AUwFRd8bMbimjLXutvOu+iXFHavfr4fkoUf5MowJKh+Jz2t5tNu3gMQrjt7NzhfAwQ8KyW
zZZmAiSsfgFRI6NhgXsRmTi7224/lnEs/w/8MksFz8i5vb4RRy9mPNSkXs/M/Hn5JbeMSaTx3RGq
rMtFRHdtTsCgYyIiiLn7yxS07umWfVORf3YD1MRtd3q8JjFAN0yWyyWFG/f18Bnxn562abiuXA+5
YX9iNxRCGBRy6LznQJYizyNDkSRU+kOiIcUu6dTEHxlZMPM68vXZtZAmI5EDLfpO7uAwYT6cEQde
sZxS9ORuFuVtUnwfh9UYbxDeNImInfhghWVQ0zmTg4+hZ39xptXo4EWcpOTQTAoscGVdixuLqOFc
GbFXPh5gmTd0Q4OxKitvCCneMd5Yu4crJd8cld9MULGNGc5d5rXwaFEOpvJ/s7AP+bOmDyiyCJqz
tBu+C8Vpiu0gHn0RGwUSlc+oJr8RTbl9b0Ln5MP8Qt2PhYjZ9/JDsKZy9YqFH/k7msEZEhKYThON
iSX9In87twgYIcL5dD1SBitvpoAryh8TU02He496WcoPVD47I26eUhcCgeEuHb9Mc3LlBKvkvYbx
asEqVlWnLbKlZWXNmd/c8Vd5qZVZI6UAzOlIPfv4+XFQJAxogbYzM8Id4W96lKmzf+83T54pDbn1
cUynxkvS0rUZMW9htPhJHaqdOuxXcfsAXtQkjCNVCIjMxOlCb2OV39SoJmVHTwIPqaUu38BZJkWL
apZQe6oWBX/MQOMm9XbSzWIwU2/Tp5r/9OJymK0VxQ5aBHO0Vg7i8rt3M+i1qoc5mUf7BPl4aVc1
WeuM8nPJCSUQAtja6EpcjLwNEtcP2sxOQSBB26E2yXrS9qcn1LaaBGJKBSVBhH2HTCQ+rsvEALcv
hAyyKhfiKJW0bABSm0X2H8sv+VcS9pJzP4Qvij8XUuehYn8mXrcuoJ5Co8/WH/bLAIIrf25h5OEf
Y9MKQkPUu/XJnHj7KAMqCqWzTpQMBa10z/8CIWoKf06Uqs0zdnVO/lteAqL0HeczRRTvboqDUQAd
7ZMwhbPMIuxp1iVnTegiRAfpYvBe0GAi3BMCBrKuNDYKrVdXQ484q2YFvnIK5chwL/rkF3/tuDXz
/PBGiiV/68jSxjTrodkSaKwuezn3Yejd9mJPtzLM/ZHMWm7S889HPvamulKBjAfSuLIOecR288dJ
d1cH1jKMb1xotA8yWHHKU0vwq1mINFWwfxo6azvImhkyYZCvrdUvXzQEV+zdPbT16/rT8LDrCLid
S9OYv6l/Ft+qVa5426PsvcjscShZtAIfKXwNaZadP8V2kMkmCGldgtdhk/ZTk59+RzKxoJaDGjPI
A98CcPGMc3ppvAfwXbp3r/3e7mHg2Zox82sAf/weYnff26YPgIOCc1LZuVP4t6KtU4X/xV20ni5f
4+tJMl4fUB2pme0/fe5CXO8twN+/ANpcpORL6747Q5AbGIkV7j1f+x/R0zr0dvXcd/5IF9g6p8up
zIf1x21tx1JPxgAWoN+N648yhsrq0rTKL0YMf/xsNAgjwxQlYi6hBdJrJvvR7zr19F0AkbObDppK
BtOIBf1NblaR3hfcsoResjcJiu6znPVKxVk8eH+poqibL6MA5Aa0b6si32+lWXlVTvPewCnHG0yf
K2mpHM9OsRtIUZ2/zve0POiCeOxZf3ZS8ds86osNi5f1qFNF2CVHN3mzcq0lTpGZbDfmIi2/VveC
nULieLBRB6ZYDVeAT2CGDCNqMnFlzEY+BIYKXoXwBKkDWPKKr4tobzlTtQAdfpPWjAypiG7EyuZg
UbSG593PWbWXDKE/IYmaWP8TRU8GbnrOx75+3ArPfBSND62YI7trmFhvzK2n89PPyWgtUwV/dq7Z
j5jgMfn3wyvjciKalaL9E2pgiCKYxWVBEu4lMnSJ9MzzGCVoUJ1RPteRFmzd9qjgCnJ7q9nguL5N
o5gtsFafup2NHrTlGuxyPlcRix2uy8f5HDuV+bwmu8k7ZaBpB0Q9kxq1tzPqiRMCmwZcC66AXRmD
SeNqCfGezAtegTI5txDUaKMPoEWri9+mEa0Dy7rBnsArcBaXf6RgdX/4Ub4ec1z03x4AhJ3JJ4Ea
27f5f3HPvUwyC5hQd8k9dT8Dd87FVgl7iJI2QgJcBk/03jiDRq9dgpHA1owVR56dNORF6Zw6dAaV
KF6H9av2F6B+HLodYUV5dDL5qP8cfuyH0fjyztTWx4xDbMMCTwBLm7i9Lz+JF8DxMuDGOzAaYuAU
n1nUNxfXxqOC+IYpn7I3btHcxoaEqZ4tJOh2Ys27DHhvrYDldcrnA5G+RLsiGMLbU9l0nDNaVQhA
Y7Fe6GJLKRnfw3f9OuoQu9gfz6ValblMBXGsl+ndsyRNi3tEsfSTT20bE9y3Mf6URrSsMfHUVR8U
VeAbvU8qwCYL2aSC9q3xgxzIMEH2W7fqIEqUf3eX6Xd3e/eErDzanDDvHv5egfQr/7ZVWe71WK47
pFNFpuPwY2f9E6Qu9C+ymrVBwF9awc5Nq0zuMd+cI1k4sq1nH2aXAg5vqB50kjQiJHHDTALipvgu
52KrQfE0w/sfwhSxqqBFsErBmy3LCyB7t7AB11q42odDHoc1thHPppoweUGSNysyzjliq/JXdYTL
+hOx6lxWnc8mnT/I7UAzAUpgkwtrzNqhnxaBttRwgo47xlR3g2kT2A+G/k/MzrjzcIzqLWiIDds7
h5Xy02mCENNtHZLVvx4iy/MGBwIC/lkpBCCZgBRyofFm9501JszQtZVqSrJsM033zf/NVLKb5bvc
V126Do8EhFGbg0kifzjTph4CX8XfhkyDpt1QLlYOPlUAjftInRUtDHXMypUlyHT4Gp+io3f97Yd7
hmVf194xvUJbY7dx3dfyyUazHrJGgsKG8KsgyIeB4QZoRML/xyk3ua0m/Ttj0iaRS98GuHWAZPlp
PCb/jPDHKxTtxSAnSzAeXs4X2SoszdbtrKVAXT89r1mPQkuuZHMuatmt/3MTJTdGPyN+dpta1lv7
KFnVopDKCRcQnbngxtLFitE2GJ16cqEh3A03Z45/N/+bLeqWcudenlb2Tieh5jGh2/IMtVTZLkLU
VHeNbCLGjD+J9X23i0mZDu2hz6Sb23dJJMXUD33LB5SIvkiI6yiJSeRZnlNwOWqWEowIQDZ3eYv+
CT4fcz0X3jw7OmH/yoq9UrMo9uGsywIApozShFMzSkUjFKdKSfDWeTn/hSyY23bJAWAU1HeYbGmZ
X4E/I6lR0smKcTQ6FjLNhOZ1DJ1Jw8xUBayMUsIuo6h8gETWuDWY6fQCOKM1M5jaGP8np5V6aF3i
9+XIC3QelvtGX8CZKri7LHmV2hBw7nsiLaaObI3u6UT11FReqLrpiMKsnCSRdYKDkse+pG9cM9GQ
yk0xCUYUzOhUiW1n1c6Cu7FGNfoIg7lIzhCka4Xf+N2EzJnfh5zmEjMIWi6CCdQA1QzGZ3EwF4AP
ousR0Fm2YoZmwbG9lMvVjkTx/sSSDhZP86Sw463k/Op6tC5tvCtgPieJD+GnF4OtIlC0CFJoasxg
M6rBc38iLPg9NO1SxDOSD2V64AwT7PtYWVlQF41b5qY4ope3lmbL+z2S4j6+m9PogDTKFF8DaBJv
hgxK1lnXppXIwdNnzY464C0q4nTQQzbU8uHQ3s//H8ApiAV+/iKP32wD9YPVGvYqzCKKOzjM+eUP
Fv31jVZkd3pPK5PqzOwMTLdGI6eP/qiUk/cM1fb6QtFNtjGVC6ptLD1mCs98tqnCHyLLBDkotx1S
lhc5uJ7Jc4Y8WMohe3/dWr0b0rAis474cUVtl/s9PVjD477WO8m8Ddr2DFJNgwesg2Jcm8yZgNHl
nNGvUiTL6NQdKsg0FCag3rfaQeURlhD1DsWwv54xtg5S65xDdCiQRHjqzfcdrs785IgyE9ob/QGm
hqCJtcHYhERMuNkiYIBq56KXDrIJW6K8Lx1PMD7uC/anpJ7GJtz893wPJPQYMIWcpAq44gGkWq22
jxibF5/KFaIKMh4+wWpmygxh02KCMjvE+621d4tS9oVlefHf8wY6jPLJoMVBbHRCSKED6Zfjco/G
M9FTCB0rTS/Zp09TyXh6pU9C7+AiY/DYBP1Vhxc7I1Pz8+HAJvt0Rb7lL6/8JxNFaPz5PLovxgTN
VY9YPDga7ww1E0ezCniO/8QzcC5MT8YsA9KCVx8f6EIOm12cpHCrzVLUS6RL3ezS6Jsmg2xzI2qD
H9RCmDA2ASgmthXdhuObFUZfmJs2F/0s9uC6ZMMpcc0/Cx/jXr8ZMsGhTlydHUH6ofKvKntuhd5P
eSneVvqd/rfJh5qAq2fNwa4AYPmsDllFAegezIxCyt+gzizJScvpuIxnIyuDcdbkPOHwBGZTf/ug
xVEIrr8g43Sdg4I592LqcuvPAhX0tindF2y5GJKzPy4iEl0fFXpLEo3UXa8X18r06+2mrh6kQ0GT
VDrI2HMzl0zYIGlmzAfol7+2lMbwZOIc1Ebr0g+qrXfhsgOQ9QYGt5F0yHL8Lo5kDgfW4isYJCDi
Yy/onPJfDn82FG+ueVMcUNhST12weUoUX9z1ZOH4qcjtMHkEnF4C5WI/tIPuURLG32raGgEwctOo
OeX2ngcivVnyW/dXxyfsLsImv2cdjeiKgehP6a/h/tuh9tkO4sPxxX8rHunFqSP4ct+N1I+PtF4Q
Qr1wZJA9w3N/6EUlOqC/EgQM5UDe9d8dk1hCYsgAwtiT89vnyv/8tgCYK1bxcHoFT2YScLpmTMQ4
ddApjiB/Pz5CMbzyj9Zls2ryVsfE7eazdNpW/FL/ZC9aZFLtGHM0vfmA7ecxqS6sC+0IMwtzF3DK
VB461jSu/TbqP+3qO2gBm1qzNPEkqX3WLsXIeGN8qPwRlIDc9HCfKaKbtII0r4z5z+UjXeKkx2vz
t6ZzjSCiQw+eqswN0JkYIEGTiQOlYHvd60kmSy0p0jz2KekdM2XcvT62w+vTR/83Ni1x2VDTOyA1
f+5AWUEeWmuMgCOwjybbXSIhS4U5VqodoeX7dkqaoIK1jZrRaf0F7EWQ7ZvtmzoFpmKwnrRDbg8N
8gxnvnznX1c7jPKpPtByfLqiFNt0pYv0m918H7+3Cb0mfp5kYI4VP52XCTPsV9M8RYesD+rzkf2m
FLsdMmICH8Gvi83ebfZafwXodz03jqWkyKshDtjPrnYPErdf7hOQ9nMOLfHizqC9q6akIwaSi5V0
9LYkZ1eY/K6iftU/e5avK8ZtpoWyEJ+pzF7xtvArojQ1t+Kt6vJJ6SKh2pqPQkN4BtUDUz0Y4nRT
zmkWTFlNDh0dhriSgatMQQrR7O346rkN1JaSJjrKy3GSPKeA7BAYmBr0YqUEb8C9TCNC0q5iGWDC
aoV+/UQGZhMNXJ5Wed8srEM/TrWfKbPBk4qc9gn1UBopfUjv4w8Foa9aF4KgdqaY3ng0rs+o+Grp
slGWVF00nUBhDFZc+0524iPhYuDMQ1wOi9Vwcy3acoWFZ2XNlrs7t540aBLYEEUq5nFZJSAoL4Ko
e0MrPU30rieiRCQhqUsCv9dgx5DavI4JAX0wHGDxcZRjoVFRhTMI/hFRGlbfps9DpIEu5ctEHbuf
R5J6HqVXSanNA5KpZGneHpXJWo+1tyGdmGPow+m7cZveMrjf4TLuJtN5F4GyaNJk7J2P5MhQ7y2H
qdPP7Th8njitADp/SLjL0Nniqq9ONXMfozZYePL7FGlvj9fpzJGoG2ecwH2cw/q7DKgiT3meKa4r
cTCGk46rkZeRKegxHNtUY+9xoF0/6d3Kfl41VE/3t0w6kVP/LQrOgDVwp9fP29TqaA1xSpi9+hCN
6UVriuSZUKUoJs/lwPqj73aIChNoJJL2p5L4OO+oBtg3+z6Aczu3JLpNRXyztNIkhalhpMx/4SIJ
jCeqaRGxXx0JZWnuuzxIzhwZBZ/I/Lk8mxBcEoUf+VfKqxZEMbsdD/zsIHg+Ex/GxyS7jyF2KB/3
os0vIch42/e/N9AJKnIAVxAuOf12J67ryiWBol7BDOU+7QykTM0w6VpdVbQKsWsIqO7TnwUNT9HP
iJeipXV7+U+3BTtZ6va0Cas9DxSm25SS/q+sJ/MpVNHTe3JCBRplIeRNfp1mSozsP/hmHZJvkCBY
yt/Hos6/Kf6fUIm4ob3yr/InqMO6HH0G9veeozy4Y7f4b+HKBMTvEvAIKvhAAIGWZCwG/8Cm+A/q
OuJoYCyvWZtX0QZSig83HU6JfAci0YOump90iCPI35zBoAYACBRNqpN0G2p/p1kh7wCt6xkb2upn
ymMDo4tQu1ixiEm9OY86PEykiYm1eeo8Logi6qE6bNJCc69Ucz0rZ1udUFKK6SH0nnPuUjJhyCHG
OP9SSWiki7+LmtmxIKCpn9S0YhlSNKlAeA+1I4Zs9Kun5Ev63Y8NWs3VKtZl6ahuBVN7wGd1HFaO
Fk7zUlx3WzJLpseH4smVhPcu2ht5puG/nM/bUo0vlqDsXCBsdls+U113Zfrdw2RSKou/FZSKSFd6
3x6lRFwW1RGrRweTtWhryEexeao7l7AWobBEmtsZ/yUjocKB1a1HJa+RcXB9iLHmxyHJu+jbYBBo
pTaslYfXiIDWguwXU/rnMhNvJnON8XwlZ61skxTPwcsl5ell6w57ylVU7vUL7OdIMkg0Gw045P4s
q2T9zj+qG04FptEXfeG7mj+/nJA8iklOjXMVPfmRlqoJdY25mvW/aXHTLna7eBCRhj2Lp92bz/Rh
fkS4c1m7QksiXf0IAtAkvy0TmbzX/h705OBYXGLKq1b1Wv/IhuyvlCiHe+JAAm8v8FCk5Fz9mGKl
LadjB0hfKYv86Z1ELIZFZhzrukYx+kjfWIkqE5ULDVDcO8jYSLVUUJ3ihPvctfG6ueMsX1Qj0bZl
NI+61k6ay/07O/Dx8o7WkhvbV1nnGHHTfiDpx5GcyW/Yu9322aAur5JVxadrhAKoKwOKUXy6F+Mn
LGQZI2Qvca+9D9MOl5fN3ocyaG/+KaPYmVDclFg+s4q3S/QMZiK4ewnmpq6s+QksoG0yegyjwW2P
hrZ7pnc03vouHehdrxWvcGx5GJSX8j/XgrZwTsdggIwETwSp1k7adNveZnTfb1JUCOliwqm9lKAy
Dn9zVkmgw57a2Eq/ZFvJdoy0iLMv8W09dtZxW/wVwsSnszQiXp9OPzcKTELAnZv7rFr6bT+JBxPy
5Wzbv6HT5mznjWGKpdazxaUzJi114alpcrn8v8zjQJeZPr5mL5QtfoW4XdxDGpurNg+3DjwPey6W
NPf151HGZNooyRuMGNwSeNJ+DsaX5OV4+JXjN3r9TviRsXNU1P/zt92gFKSkeAhEk1Xb9wW1WY37
DoeOoK5MCozQC84Bc5r4yEHRQt9UKGhkur852EFIRaTqyp3J4yLkyOpxtPQicX1fvx/efj/wxxLd
7ppDstHyPW6YJwzai12neGSF4OGoSu5lwro3+izS5gi41JYAnizTYceAw9FDGQOcNGVWoIxyr6ht
vSWtbrEhODWN0XUezYzupTRTmuLPXrr2aq74xBRQ08GdchPIYt21ImkNufAjfhq+oxOyAEs5ixOD
6hzQf0IRMrTsEKPWgrHNFk4tmPoLPG8YF6LEA2sTtJw3VZg70fRiHlKztEbaZA649nmjIIGgP/Dw
G0IQSm9CpCKTgek0rUjew9eVlsp06w946f/C3ztfk/ZLMXvUOdwI4QpldJ2igZKrRfr4B0UMkP8O
N5tlAregHJtFS4NnJXL0SlJ/BiMaiOGJagyh/otDc7VgiSLR21olhWZisOEI2KaOOfS5rKw5VYMN
/75obKA0xXU+Ins9rp26iDF/eEJPVrpz9znm6PmP34ieTGUTn376PHAkjqbE85w72JGfp5zzAT8L
s3+YrcE9GEhQK8EF73LrAu4UcMaBuqDYZSiaOoLfaZcPw6xAqDtoAtM+N+JW9AOTRL6Dud/lyDBa
+l0JxaxR8qCRkTMyQP1E6axIP/vfH+0SGaC89UEGKj9nM8bOejh7Y6ggOOaRw5FnBUIYLavVQM+z
xxKEoMpn3pF5+GN1PLd3uoKtgnaNKX/nhq8reNe1gjpeWH2j8xTqbeyUtE378ibZv2peA+57BoyQ
g1iM8clCS629mGMYsMQkv/DOiGCgF0fc0Bp5+8YlGwPY+kJJwRvgVCIb4jG4pjwaYgvfiE9aCcr3
bq5svsc5a/KxxjpUEQpU1VKv03sG4jAHpLG5YZrP6GGW5bxeag0jggLaFAKTAoZvXBrdlW64/Isx
Ai2yEDUty/wfXo7H8IgJk7BYrBJY+ohi4JoO/R7zcKsMamtQGnQAGSjpq7g/ftOPIUhjCMrqKwPA
Orl7vEwIq3hPufkhChCVGk8zDCLPdCKatUaJ2dnug+wHAZDC86ncRl5zSCWIEXS++sMqlLP3f24L
Tc4bZVcW1vuc3qtaQKCm3BCsjqHCR4yHhkVPSfFKabdWOWvOPyqGugdU7vjQvXWu+Uymzc7AhW8b
2+JMfNI+UU7kW48/lWcP/njdjLyPAEAHq2sJEdPrNG0VevuMtcVZloBn5ObamOkQ/3Cog+LEXsL0
Fp7D1hWk82PZywqcRTv+gBy5bm4Y/1Imal0f85iChzffiyawOa8zEAHo9CoDQPbNw9EjAzNDXLns
7Y9WfHcDVlQC93spBKVedEbYXDmc9TtVuVni/jNguaBBs/zObzB1QYpIT5KakfRZmivk3lGkYgnU
09gEnI77cpeTXAfubqFklLEmoCF9YzHSA0JPbF9FYQdWegINvuNqcfI+EI4iR/8rNg4PVCsMKJ3D
ZpD/OwjW4gushItm4sol6jnVlssCIwDlZvPzL8AXirEMv+nuKvH+BapuIdk60nA30Gfg3a/OJksk
/UUKgj1ujpYDOlyqT8mZWm6godzGtPzlItGLkDKPnhBV87T9D029L7Us0dct/ealoc74Ua2E3rTm
Mit4RlzPQPbZL31vPGEkKvrV3+F549r9HRQ0WnBx1kz0V0Mgrk3AVZ0Jag+uEEEXUh8mtmbs1lcT
6IcZSMIyq4b3r88H+EAHmphbgrwtvaXIiCQ/WLE1qcDy5Y6idjc3pEARuszWyF0oGj3yfdDLFdnf
1ipxJFpzc1+nj+uNQvEsCLgWkQ1cC5W83+6pT8wygjI889YYE/UehZytJz+OfXLfYhv26YCai6Gs
KSu8dEOIuFFVJgyBVrcfG70jGM8Qjz+lGm7OT/SWCFDVgMROok5QpyRmJ+Yd1BtzW9yWOZ6Acsq/
AnJHotphbt1o8iMp7Q45HkJq9AdEFTbz2O9gRU68SQ7dYez1ub4HWbqbIOb/WDG1r2R4L8XPOWO9
AR2XiL+BQeCA7I1THHmUdkJf4ef1dnnSCEt/kz99rHU3gW2Oq52ByZiNxpOWX0Bci9ftfZxpl7hV
iuYgq6Q6Q3qEj4L1Ygf9gYke9iQQbF19Okv2SLOXXwo7mH4YfYdEmS5sD9hXqJ/wltPioxdzKd00
9rDKhKGKJGXwgLgomszkR/XXQwlZTBJ2KRDsXnm4vA83b3biehmBgE5VCdTT+HWjdcbFKLnsLR5e
eOle8wQHNSFe9j93ItmQ9U/Dnae5SzqkKnt9u0BeKT32s+ulwrxtneT0to/T2g3Xa3hHe8ol2enf
PjG9ia3byWbglwlc5cdaVIG9DtBsMz/6aFGnVkkumTVoa5kPxmupe8p5p981A3Gm6e0NGj/8BCyc
CPEyqNEdGbxDSrZtqgbO/v4ubicNqFMjnlOhrZP5OixFkJLFZ1+6iEIN9fIPF8eDPFnocJXhdU2I
QFuXc6OztrgmbKITZfTm9N1ujGPY46j2umbQ+6mHl1DpuOrn0+iBbfAM/I10zDyQH8KCzW2w+8bd
FGeDsu3IBRHtsudFhoi68p0zt5auoHh+Sku5H/t1W12IJZ84wKCpUp39rVkHIk35lwjGjb27rflD
K1LRnH1l28NNP/rPoYrDimNf7PyLskcTYz4JQ62In0M/O2dlLdllYY9K6fv96jkesMbWJC5xcK4C
K+hwXOpEmQYQrAt+877aBGNmsMFrQg9D/Iqz7Hbmm1sLe642BF3opFKJExPM/f80dSDYVTgftkcd
rPYn4GctZydJSgIhIZmKtUx6JPqbIR4a1UE6sXdxEppTySAEM2NUKMK9fwuRCuLMtazXZTq63BTG
ExIUDZ4KbYq9CVsibf623W8Bs9DM4fGNMA6vZlPio/CXJwTCMSB9IkZL5/5QeLZW1PKQpPMub+ox
purCPG/XDCXoJW3h0xfB+0YXWk4/JAPnx/G5gVTBCdzz3eQQJ3xwA4OgWCFEq+Pc/OC9knX6fq8P
f/4fvPFC/di+xMvVfwPhOKrKQThrRcTlFwUU233lU3o3xxM3x59a/ngv1N1uF3Bv1DZT6FkrOCfq
vh5l2TZLa1L48h2wN/tiNSfZSfwsZnZVH0Dk8rjJ/NECcPiwLD1UU4TzsnTAfdwAUJUJzq3mD2oA
FLT3+OhgmhK5ajhyCH8jCTRkTgUE1MvYtCeyTqv3PEu1xcUO7rfkYLEp2MFOjHgrc75MPPOx7AkC
NiV+Q1mWg5ZHM17m3Z5YdWQNdgsa4plUOBivFHQaD+OZX+fr+iaBLW6CjU/UFfRpZtAoz0uoUZu2
8OjGm7oEUkalkrQUYVav6EYN4KvTx7i0BDxt6LqGHMX2Y6s0wizxbY5cUSBg6tTmkMpo5S0fuTse
gJbujwzv9A8z8pslmmPqDRTeR5fd+dxpE0m11GGzeSJl+6GpN6sUu0hXbQ/l9hUCP6j0VguH/SWc
SXZcLYIzxPLLPMqKLlN9utqcccJRxWrYKYPAfTnbapfvv3DK0LsYtO3hQ79mSSNi5dF1wftWi8/H
Qt16fdOqRsRuU1SoUPtTUi7LzEp/Aho0yQKxqMgBrHE=
`protect end_protected
