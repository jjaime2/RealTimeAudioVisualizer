-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mqBKKrDVpCMHWPYDCpQ7CgSL+hzR6R/0648q6BCFUhT5xtOwtjig6HLxfkqp+AbswktO/JBrqWIA
SW/XIWXSvE8+EwuRS+1frziZBk2x8G1X2DITfMgZxFFG8QgE6LfiGAQWIjaafg9/rsgpeylfNF9g
fnS/oMobmCbzomLcv4cxsvgUcdQMJW++XOIxAKoEptQjVV0kOiRhwsEulM6wAe1xrOdgVI95pxif
TKaMv7OWMdR5UQBY7wmc6Sqn36BvCuujwaScSWxgazF0fHeJXxcaqqCC5L1PNkLcOlthl3nGPF5u
gj4ZPTms9pcI0XQO4Iady33IWZ5tkuVIqqnZIw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9552)
`protect data_block
BQmT16WALtJc7emMUaQmEXx2Ei+zaQmf7OzRtICsyL+QgmwajqhvbcyuZyqezAN6lipqG0/Ds/mk
zCkEG9xbpl6maMB0BGQWcniJhhMf1q103xG/8QYDjDKLEu3KQ5D/3bJog95BiSQ0kd3vLKuDjNVF
7ZXJTP1+dF5eTsLXcxc+/Khbw9XCz7vVhbq6SCcfDHCmXK6fq6O/Yr1kSM5/3/8P4L4O8R513tO/
CMRNkJ7Q/rbf5Vfu+Ta/0WYTemx4rtwk1L0Y3AogZc8aAlY2bLXeRkluW/j8s9EnlcmdjcKQWiee
ulK1ixelWg9dkhtCD43Hb1ffFoh2FqwZeT+hFFyhZQIoJT9sjdVFepu9ogu2Xq6BLXGJqfOIfPg4
5QHbelzANRJ/sNoZymkzHfIE/kTddqZIM8qNyRKAza0ukA5CxNaHHH7qitXd1y0sYWkJyza9QVk+
eXNtBe7SUSBWZ8e6V176yWXbX8hLEcoGFLo9EfQW/GyGC3phGB6CEihxhR4Mbmkfj1f8b6GXaRTy
tLljAmKum/CZf6KnL9JuWXQD76qHkcm6ivaT0kL6kJt6mjp8ccj30bGJ7UoAddUnu825MGjSJEvw
1u/zpVCt52QlIRz4RG+q3gACjKRmFkjB4ccQrwUkAF71RGt5cS45OvaX2UI0Nd00idqn+hiHr8FY
20njLqJgUPdbwRxFHMOugXbKMwTrtcse46Z2gnFm2tkpvJYBsBx/ezjwM1trJJWI7liWzfajN4Cd
W486zlP+YwoB5/Bzu9j5yg4V+P8goIuoVBgoUgpYHPQ7ppCqwSVAAaEmOUuFOZWEJjaj859vwo3Q
AN7CA63KTh9B8qrppRDsUvpM9pnVE0lBTed8u17U1eLuNYg7JgXI8O8MdnX2Xgyop40VZtbCQ1V9
naEzeb6Khioh+ISBxzsddVdCX4KeRc9La09zgJ+yO2R1CuoocgidndBkkGL+E9JSMUOJpPW6udZG
brc5wMXTQT4lzEYeQfzdOqTlMCHpZze0IpAJWy2tXIW5+8LD0hBfGa8emJYaqkCUpz1HkjqY5HHr
rJTsVvbmAgEoWSz1RnSH3sOk5heTvR/Q9pKZ/W3sJVZzK5sUVH9glVgVXJqfTksQCR3q/V7x958w
ThYxMrUjvvMPrSOTdMdrGQGW9Yy6CGqvKu932M9HNpJ8bJqqmNPkdKbRp78d96FlauNbZz3YlpdK
G8V57RfEmzZfkmAaun5vETS1tE/ZxOB/TccTxUmWzECB0v2a0jpLM0ySexcLA+TRYWvby8cpEDLU
Js/t6mq6wR6EHZ7Fk5Nz5bfazXGcbh2jpGHJ/jjHZEVCCLIBAp1kAJeKjaIIgeW7sxrXkNOOJgdq
2BxIGLwov5unCzJtYS/B5iWfsMqv8Bs9oo4/DcxTGkasw9DQKd0jpGPmVk1aEKuSIgZk+aNfJKVn
wJ0Lutk72qvt0/oBhbZOLUqpthjUghDthh46eH3CQF+yTF6fQiMbR8ue9tuys38CD6OGGinAdoNl
szQBFCIv6W951vMGXrM/VPQo6RBA4bIMnoFXDzSv+wcbne3rJCgga6bL4Wu18sqDUwqTQswxWnPg
3GZlYHRNKmrpvn725+k6wFhhVcYYEkkY0Ytz9dORBI4lNsMb03nulvMKNA1o/K293wm/aDWu3E73
0olWD0FafFMGi8OrSzjgrX/MIDzyu6Sw+XIbqJy8JQ7TZ58krMZ5cM7I21QHZyBvPiRXHziNNE61
iRezmQ6Z/dHZaiMngCSHuhEljcbqehDHRWOF+gnwI3z4sSRqQZWKTckEEMJ6UU2w2o7OvN6OKGmU
DBMPXVmwpByMqmdLxw5rPzhWKL3Wv0PoAw9gVYNjZRZrWw43Bn5UG5k2aTgkQGQUMaAJRyRm+UOn
BmyFkXDo7j26Uk6Dk6yh7a2wlLlNR0v4qAHoNI8vFCxvMdoWM0w67bTeGveTZukO32fmID+SAzXH
gb0LkXIbSuu5ClvDRpjd6QQUHRC6xIcvRlSyv75dQRxkjZosJkvotet8fhY/lmCpoLJT/3F8zdQq
ymrMBHgh4wdjO1c10tiWM294QkjyXQKgiySQbRb0fFi6dA7xS6PipLxilj4VPUcY+D+cAZYxOmxU
czt2btPZyxOOXGrs9nWMkkl0be8C1uPpOaq9vHAo2mxDQ02K1E+uPQ6xrHEgnHIBROTPL8XlySYe
ZY/WsRm5aBRnaJhKj38rk7ob+bO8Bu40AciN0HNLCL3QuPlR2WLb8B2OwlN+Y3Z+5SdPRPMakf6z
JUiL+Zyncx2lHGGs2psADSVeHiTstM7MfOmvbQS0gH6mNdyjQQw8i44ADLxYZPIL6EjLOd8qc4cz
DP2I1O8ATCyF9MsxJZDxS7IxNMmmAWOJoeFNhn2ZdtK+8x0Xy50lL0xVhQdCbFlGb+o8nZpw0BiQ
P4FGzY60W8hLMZSstcBfF1JnF9J0ENOZvCHOUZOLoz8tFPP7wgMqjuk33PerAXRVQo1C9wgXlK9s
WwUa6y+o/fr2RsrbIrYFCr3VnqHJ8tJXQFBO6YwWKm4dK1N9+rBy3tDWhBqUs0frzHvlvqBwEI28
tlGYrlh45tFE69byjc00iuV4/z6zt8wFyfCsSdwh/tVNJdK+9Hj4Tjsio9T6rWJaHOyM4UzTl+ba
SFuTPmRYXWqLkqrQJ3D+ffyDBmPLRp1qpeyYLs/SNVT1r4tsomKaC533k1usZ0wkqcP8Z89LyJOH
3RekftMeei2HwneslAYCdpY5DsFg3fGENB0Hpoj5rKyMhvjZmu71+9R1lSxq1QH62828ZWKhQVZ/
rTi5Kcf5++wtDLW0yixzcHftEIPL8BW0v+h6B7fcdQ0S+XDDTfhO/VR4NgkaVzJyASJWzMCxq9Ta
68gv5isJb7hJxQ3LTYtsV1TBD9iHbP9DLYllIbig40rhKBPC2cD5C/S8zSOEPMoEEQqR4pIfspe8
Em/QjgmXtvL+oGUCuxCdsq6ok/iJghgwmbUDAYI7fYK3fK0Q1s+VvBpm8EOk9Fc2/LPX+gHBWHNn
u5Ri7mLZXrEu47OA1Snohj8FDoGSIa3B55wOnByvayPW9V7ocEVVolFBiEwXTvXT5NrsqYvcRGy8
PJw2H/F63abL0TPWnwJrjPIsp7EgkxmyyfiLIzImmLLRgRijIj3mYshzdFyhK2NoWytHr85FsKOS
I8y/jh6HfJIiDsx3QUrkqNVnctzli/O2OQ+BcsyYLwkfvaI/HPEM2X/kpecSZPZmpzsiVEPdLdke
8yvbUROSsGKmLlByw3MsX0Urp13V89FHkuBUZ2kRPodDxj1+LaMP/lqIk7mEGX766EQ7mI3XHokt
ngKYSKdyx5njyyGAjmbhWTD7vkrkAa1a4sfp9iFVwouQkMdUUd+lhvvqwfh4pO0kena8LOjMLlQs
55AqEHlZtfJyQCKt6rVfbeXyJV9xD+/+RbqZ3bup9KKLRnuvUQ926e2GGNg8jtrTFMDS7WU9bozS
FbZsynjtk6PRSykGcKQQmkxS9sALGjHV60zvZsABZYytpmUI1opj0U+QnfRlEDdu7HFrHlCqQJQo
4IVed+ypeawphEyxSixrl2wCYz2O8F8yA1qDLvXB/BmDhv/A4GOMvHCyXcoy0luXLQFWXocRgXpu
dFdo4wlijZ0ETMSoK/7GM9NJ/f+OaaR4MkjdUz8ip3uyLNllUQq3Ot11z/oYqJVBpcbOvMYCsLD8
X3UNiTuuyHaN8/XxYc7sbzmvwNJtxWml1IN+kHNc5XScWJWmOOyTCzJGH6MDtSv+svmugBdjMDuU
KscXZ/soeD2ZQj3zMCH1E2ZdSzj4/hzGNNPcMquFduE3h4AFEBSL1yi7LOaU6kzKqzTSPSw/EgWV
Y3vHddVrDJcvUXfs8cZ2ukXkoEvOAW8TeZL0mJikSLSrn5NHJS7xKIDFkUKW89JtOnFtX97rB1Yw
njHk51bfnDWfLGOun4PF3NC9PfnXx9h1Ly0nDl+nw4tW9Ew8gUatVy28Bqscf8GLHael08SbPVfG
2Zv1wpOjmzK/R3jMt2jBLLXDn8S4D1BkeYb38M8VvNd5WpZFtN78bGNZIJkwwSHK6u65lO+UGoq3
PL+Xkp1PL72/UHyQ0pNeA0/IAR4i8kuGVi2pBFYqx3IasHEJIcr7npIiZWnS8Mu5cvjTdy9EfnKg
QUqbaH3t2iHPD9cAsRg8iI8lCLYMQjV7rmC/v6Qwg8ly4pCi7ahGma380Tiym/EjBpHwfkPAGU7c
ULhhPjiwO1/JEmim/FNbyaYlhaPRkXl5rbPW5M7Hc3ZlP5qrpJeHA/o7O43zVmOiRf6ei+xY1lH7
IxYLlOUD0HIdkhLBUsttMxVvF8Cr9RpivBbYw7XxwD8cJKLljkzaizWul902JXQrbTFrPw/lypy/
WrIwZOybvo4aRGxcsVk05LiB4+jjdTcP3M+H2wVEGsM/iQfj6lSWvidf2HwVUtX1LuEydSij2dXu
Yvfl14Vyr6UGXR3TFhsrRx/bdXKKyjtZngysxrjSYdC5IJeeolmPlBgYlWqW3FY4j0eeYafNaYAn
3ecElmZiUS5xakYw6FM7joJEy+8xyeIWXylEPSY+ztdvrEW6SU78QETeRgozhAOPHi5ghGvdkNJF
ZHFp0rdO+0rr1vghwaRSwsPEv/VBmzr8WdfK+bsEfyWMaYESLFD/LUUFaix239eMzykWFJ2CvAaY
PHFRD2DweowxYl+On0xXwv0IEwXPw2b+m9guFrvHtmtcZOgA6CRLSifpAz2klf8vlIbxjOh02zi+
RhPhb0lCvK3LjXJ2iX7T8uXSePHpQUnUug3HRa1nteQ50U3OO5XBpkO2T02E7JDVfNfNWpluImaU
gDjCDDqfx/eEDM7ka964QTlysFFrrknHI90fXy9ZEr898KS4aCDJNgy7i6jXDYVIxwg8KgmR86hc
KQlpYHVcvCJWHpzQtyY6e1oJMGgk3Fy+bYYblmC7QVddBJUHePx6c5+pps0xDutm+g1qf4s+xQgm
2Zp8FnYZaLyt8XKQuWIlEknRnnvNaMFfL/SPM1/RO9uTaNPuNfSasFbzULqCz7gz5zpnQYDsfI11
Lsb0y4985M3x6rY8ctU8im6htHh/rECZYo9UvSolrzFuciia4bzn0/2kINSrSUVxyJ7vCLvF6YbL
ebHDn/kUCAAazBEGrbaCvkx3QFB0xOdGA0rnfup28wPUMiIQx1BAVmSM+mNgX4AgTXrvOCMFnxK/
enFx1ubNYWylVvRZYeOS5aB+je0M8HXchF0m7ISUxnimBUbNqtQx5Iiqg7qp4XSWP4NkRZFYciKM
J80APOFYceWwHFkZ5M0BP77gk35JjaYiwtfRl0QD9LheRKjeOlCk5hg0o4fkE0YQz5czi/cfFwqM
SByNFskjG58XRMsdBfDKges6jn7/SUNnTcGL7E+6PsXkhhJ8owiv1/eILfw3th/WYSw0HRZmueT5
L/Ek9lAFVH6jI0COocIEcvcRXwC8/A5QLjlrLT/bOivs8Ub4uxlhT5ePPnLGjjgu2/+uCLrzDhHp
iHMtgM7XOjUt6IxyEvOJ9ssFHt/yX2k5dVjZ5eN7yTXiLcocuuXCpTKenuhWEYJUXKUUGgRs0ve6
k2pKbZ1+HdIvBBkaOdjg+4tUoJzdeU1G/soKR9Eu6sVY1DAkfVxjYaZX+VPSksftfJn8lFaez9wG
PuEZrYjS3nXDeawk24KUgiRPScjzNMgE8Sb+5s7mErZcLhdFkDaJssW4hOSY/xajerWotyc3dBgE
boirK7hTKt4EbF69kGeVuX7a6TSUBBR/LpeyjEKxn5sT0unJC6QGwQTyNfqvS72O8bNBxEiF1VYJ
1GDefDfczWz7M/5TN4Ne6cUSHf9U0WKZtE8LGw0oCt+B7kD7T+l4+ytarPLcTGxL9S82pUnq8PwA
g5XqE742Htjl8/gJalGA5SaB6kE+c9bQc4e3Z+UKVMFUFUHmMy4MBIH38hFue8LlHjJkU7rJD/r1
mQa1QC0arstGkAxsg03QfQd7rRaY5ohte4k7XUUv1sfgvXED6Sh2/EuO8x1aLABaKb6DlUfIv0hF
p9TdwJDGQeCR1akSAk4gVL+QBPVVeftR7AYkZzXCvAHLP+dncpoQFzGjAU53/dD4KJPdILX20N4f
Ipx2Bkk2eOGzlmEj9CNqZsCKBQDW+y8/wFSTFgsyFGLB94qpvPdXFoCbojrSIedrBY5OTsFUyQSE
lpYm9UiOBft9vgVLxqprV2XyUEO/72yvbtoAsObiAzqp96huAwuXTmKARXfJwAHfGBytUeRmWjmd
aVFnL9N4zzFfmfWBfj1dzWLG/xIqnLa/S5erQ8W1suWrtKieHBxd80bH+zHumy4HLMkdSt72QBoQ
GboiajyoMQMO3QJb3qUfxlmFgZwX3/pBwMkWyvc7L9EwqSZiRv9ea5KIvuNlcJ69sYzxYrEhcZAB
zxdU6WUBCP0+KG40t3jPr/9AdiMKtUj1P6f0FFwIZhMypRWxXXTMOqnaIrBb7dlgaGzoCpMxEpv4
HVpMIdfvGoJrYWmqxf9FQ1FndCwkPYisdbuXeDPUTPbfo0O/EGT/S+7e5wP1cYl9lyzQQTv1fRUQ
8NuQENzU/9SjF+e1X7S/PXU7jV3UvZSV4aZ9c3mK7zF8O+XIqfCl2gV/wwFh98OsLOGtz7y8XKB7
TrK9h1vS6LB+FTJ0w7bz6AxJYd5gOAjtjEbIJjWhUNiCXX4ho1kR0LdclJiMZUVX8AhzWOKgOAgQ
7FYAsjTrwPzLOzd2OYloGOWDX35ve+KdDyryqOWAtFMNELGjPcRt7f2Jx5+QSx8Rz95hDatX9tDO
LEe5n2l1AUbYuqaBlInPoCY2NNPLBlITofcbXsUHAmtLym0NpkFGXY03fcSdHFdCi/we0kkQm/CG
RUEeyVWTpBOtaFvQCKt3wAAjKf5EhcQ6fz/8SpwvAHc3yjqOhosY3xtQGSZrsPV4PofWL3GKj+mf
NBvp2GcGyZjRf7teIx+r3fM5f5eWQr/jCTx68BDLTnYy09uEZRjt7TB1LtSS+a0rRVKykVvtSYqs
oWX2ZiwzcUTxyBtxq3xY2bLyEJ3hVn3UC4bXhtVj/ukF6qNP02FlGnw626D7sbMMEaBT0TDmkl2I
c5BQDiKxfTNr7glLUw1X9SfZBI1/2Zp0xLNkO/S5uKVRcPA2I/WHonBAeMrNw+OXLcwxbC/HWcsr
ayN0sUbrZJ8DYOkSleVeJjjcgk2GCrSnmxaZpcUfJVWZ9jQoh32Qm7xH5q2MgswgCSiUUVmyt1+x
0z2GFpS3LyBVVnicjLFvQDGLgYLVmHcp9j013bqsgwBqIyj0sYVkJvwmWkTb0jMnM97JTwBVVxjC
uIa4aU9djw/6zWuWX71qROVySuyVbyHtihSZD4Hn+yhEpc86LQepX4Lv2CNd+T/tvEvC9cfq5JSY
yqN8OYqaDZviChriVhXQ3btHeOjSSo6WMyVzG6E+i2KVm2RouFNG23KsBxCdcJD9IQMw51wP6D8A
6TK7sy5mIiDGtjML23Aa9fH5n7PQb33e0wYwzBVmmlFP1vu45uYmwMYy8pNb3CWoRoHAcB9MfM8S
KldT2j35oWGKu/7ScBry8ulYxKYs3xiMfOeVRc/ijPZHMg2T0+3qogJXoY6dFBbG1dlg1ISJ2Vay
esnk95gRe3jqTXPXFi5iLm59HpIPMSPsvkPIiwUK7AuNT/ylis23bYWwv4PeplehmYeTBJQtInsk
R8JWJWZxrey27//9WhAfpEFP+xCL+mXyyB6RhfA7Tnd76Yni+zSzyocynCyvn5fA3AbqgB5dr8qx
eWRcY8cjAqm40RBLSwcFQVv1DjJns0alEfdpxD19LePt9KAdJm6Erkdeo1+4S03QKoHbtwxRtFTv
rIGGKsfBrISxRRC3OiBm65ERjUz1kkIbQJyRO2+pO2Gn8Vx8Bz2LX6i4JdCONpyl3sIEuPpD7UJF
6OSYh4RDldHEGjfSqJzzH+snczJ1LbKkudquaFQQzjB2Ocjjp2UIjwib4qfkGKC3bG8syOaBZDVM
H+0DAOk6p9A+buMlVWpdUsLJ9uNkrKNyCxfk6wtajKrOlEE/hOsvAlgaplfsr/zmbiflGe3ySMqE
ZqUxFK1gvqnGQhHKsEA4FqfnlP6nBmm1Q648JxyDZHv0d3JcddE/oMWn7jtlL9WxfMIag/CWX80Y
LstQUbODIUz0uP9ELOKJmA8wknQ5/uGv0NjcbvCGHeYSKsojP+iPd41md1liORtji7oOf5df0Pgv
EE3WQBPNlWgbKNdn/GB919O9y2dMcDBS9FyQUtcxgdJmrpu/pHAEGIF2v6wz9Oeg5fp0UeSY3500
4ZoqUvf6nt5ls5bCbkP8n1gPR5hCytDPSBm23y1NYblGlBn0CXpA3kRWwJ8jpfZuyaMz3v09YncZ
7Z9Jgpp4Wq1bOBT7nhZq+bMll/2t4Zvkt5dIly4hrI6x/Ibx4lXk0lVojnloVD7m4wqoFFDhtGfh
cPelH8GDjW0ErY7+HP/fcyQMRRhz3Gt7efh8pAbyCaYdorhGsVoThKvSlRKz9waPwgswkCd9Extc
zoDUiGg9QOx0UxKJxzZ5XoTLcWo0kHML0S3uy9LwmSzMt0sVTv8HAU5c4WMdPJRh8hgI9HxABrEf
6+fgt//WWgo4vgjNpoi22pZ9lUcGxuuhvSDaoaLZh+XZHBXz9TJabGejyo/gK6fHfftwsJB79BJX
Ax1lm7hhxTbv8ANrAGkpo2+w8Qxxli35fMgWGX9aXga4aaTYSJyIZDCHIm2+blw7MKjsKAXp1PIQ
07mNoBRb/irQiIY32hFeOZCUZUx60qDv7NV4Izq+cTr7hXMKzsGN39EeHRaNMzdYihcRgFyX1Myj
am8bQZeYqpOkpU/pYXM+MwxNkW+JmMI2jVAPwJ2k7+eh7hAMiiUxm9aIxhGSa9kUxhpOSrACd/er
8BJYFk6Okfs+dg3kIsuBUT+2xHLmfvbRLWZaoIMp6NCUkLlUNBIu/D/AtWQ/OJfxiuO/XCKhJZPj
7WOOFleHuq5NXUcpMiMY1g6KsleXMOwBy//S0oBiEuHdwEAwdCWV13/QbaHfr7/27asQGNp+bjiT
yowiQrZzJES+i6tQ2S2OeG7cWnzugAoJTT0iizXV3g0oX9zZ4rtjlw9YtCOkG5ToFeyYc8Ur5iQU
TzHsdWSfNu7tZTPMJkOCrFNawPAuXoekjuihd6rvf0dP6si7jLcBPagRH2BNDaL4xlqZHNnDe2Bw
t2PBRAllqfLaCa+gy/G7bLcmxV5kWk+n0511wHzC3TOEcrhsmHrGz+XCCa5ZMwvTUb+2julwDiNn
TpIcdxfv8q7/DPltHPWJAeyEPIxFGAJ/DTIEdPmLfsbk2vr73ps/ko/Y/btw3lthT2i9kgeosirm
dWtqmhojkBzNvVfAjzeN6FNJ8jLP3TjjOSEsLombbNQoCS4BaRXhyMg4TZZ3afzk9oMs6iIwuw6w
uz0IPb6EdfH3w/UMia3F5sl3P/eAoxX9r6TriC7YeCRERwTWMHjuoAWdlVutZzfdrrLHkml0LzNQ
l8lt4HhMBnefF9847G4JEfRf6dvQUQ5iqzzEMpCps7R86rOFTtBeddG8wyjpu5WoFPXNwjkc19ZJ
sOfthJRnUdKpCLlOZWaehe/57jxs11e5j+3vD2NbuPWMDvtzwCFJbDnxKoqu5X02O0xMfMGV/H9W
O6QGhVCWw3Q84tMkmXKf4h9psS6hzi9EhwkfFZ7Qc4+qqw92G6BUBXH9+dBdATd7iAgC0+AwimRd
IQSmrIB5aV1jtJObeUO9KDyoqJomsCfw3boocJ4XZWMfWVH30pKi4JNOvCuarVylUyTmoWjs0PX7
eeIGVBzU16yjR0LFYkzM+LIsQ3pECJqWe6ofPnqHfJAlCqnAKo1lLEDsVLz787/mib1LklyvchjU
wzhYZa0IskfK6K6wxd+V07cGBnb21LvPEEnJrN9D4u26dou8BKbTsWm26BspAAfANh6rvqhhkIh/
Zsr3CPQDb6ccfxIXsGQ2aTKcyTvFyJviqUscgCEK9WHs0HlR2PWvYlhrnvPQ2Vlr4B9EDg11rczm
MfqBh8gj57iH8hXjWuQDQWMsFdcev5kVIHsMnuE/iGXKISKvNVq+HHsaFmL+lhnrwxipIq2xeTjJ
eZZ5dBsEIAIO0jhdqamwiugBsIipsNqkFgtEYPtgKho1dPgxBZFYYeG0VKLSIWEwf1r8rHrWcZcU
yqKtXKwhlkF2GHE8SaJAJ6dxd+ezMQWYlEVaEYuW77v9QwRcNZ0LAbE2F1dLc+8C5YQFjNKUI6G/
1rQXxygL7IONlzicRseUsDKrGOSOIRaew8QNrpIXRKBKoBSnYGK/5sgPUtHZz6PO8bgeKqbOYDvV
PcdZ7gEJYuADGLYiEdSY44m3ZWp6tAouMupwjUuqYvEsMpx50JFWxk0cY3lkV3963/0uIW0ujYsy
C4GlICSvzM0yugrnlBgk0VHR7ZwtqicaG/TqnsyL8y/xqREqQ5zESwsDtuUZyB/htebCKxHRd82p
y6ZvfIAwA7HahKZ1Jx0r1w1bw/obcZbZkWGTMZv6zLanuP28T1Ne+m9TssEnfj0NafRMlBqQ51xj
AYbEQwYsMLIRWmwyTfeiWSlQiHpx5xSag06KlBuql1einiRnLLVHeRDbUf12oAgwHZeE0RHu4K1Y
L4rhT/sySBlNoWPUXphZm4EKZj5sZbwdbIT8omYa7C4dUH46mijihI/i2afYdmtaNQfXb1NBysk3
gaciZ+uL9CLYkQqBAoTskQMPmdHL0wkarpczV1zPOS/0bPb1EVqM7ZNbxzFBAiRFAVBhyq8EpEeC
yqJEUMQyyqe4Y5I9iia6nJjBGpRJ2xhms7hMEhQCnHclrtVAYK2HURBIcReo1Gsgqg6nS0HGVj2l
0P23KAnRhkOoAXlwYPLdtHelPz4yWnEQNyS8TeOJhhBGpcWxu30QuTIW53PGfu9oorKQvCzh6NIL
DERANbIUMtSm8C+wMYK+ZrLInTv4T5gnfTggKn+6Ahyqh8ZcFNtfvjplILZYOIs+4Pja8zqbBT7r
32g7x1LpMivx/KLUNERIoxhpw582cCoBintapClRPKK8KfwCYuBMIaotKw1aYog9hBawNMlcyDil
wGJ+m2cQGQ4yy8i75U9n/QY0wwaBJrib3jwwgyv+Bw8UkBvepPde3mp2iRuR9xm4iPUt3Ide36an
ggZJUIGsHQ6hk1lkBHH+BHmZ7hEcqwWp98NJbDk7z5T/0TYUMKN86DcyhNIlaDbihNbupaPyVwKu
NLw/JecUzrl8Ft9/6m0JStrq4Et0O8s4wPWli9ymzZBKfHOS6szRwd83D2AkL9oe2+Xghpuy7+Jq
zG67wL/Se2dbX1NJmt8oCin1M0XCR6WObK/vsYeMO9k75hCre3C0ou/lkVPwlUNqruwPp64wcMa4
zzkly9PuovRRmQRKG6S2fX0ZtCSgyijzaJugonKS29ypF7wdkmvvVI0hQypAi7UZTFakbNrE97Gi
6SvNfSKgE286m9DQzwNo8cxrL4VnkiehqqKrSjIszU3QfW1aggvXdZZUzT4e2RiuFO1T35ne5xQt
wh8XabvZ7PdW9FMH5CDPZEE6p2ZWJIp/VrRYspaetr/EupJIbRVTVocm/4Nx8UxKrQVmiPFiCb9w
j8RkxV7kYq/wI3LVDINSwsXSVUR+9s1xhRIn4Q/r550wjDXU5UGpdwN+vv30IJYB6kWBQJwmM36F
aExd0XC3PVIb2evU3u/5Xq2I88Ke43s9y3HnMD1JKP/m93iINRsJJ+IQaJjy4mLp6B6kL+wqCMQ2
LQlIoWE399sKVMxLbQu7+kgFcboH7UkPvUkoZ47JV5aLpXdjohjEXq6/gj7osIHCfAhGfrzYQfKk
OWubxhYJpQMXZBxVNPjol5OX58ajDEODhh0DfDUT7f8JOjl18qb7sqLJXthoj15czNMhNF8v2aAs
xmEX6ZGstRpukU92DGQMyecjGpsXx8lL+Ux+GKqkkHAX/LmDrTsx/HLjNYhbWeBJ9A9/Y/ozQOfW
lSHNxufKnPpMJrbitDvgEhDY+Q43bFH8c0fx9V1pGSzqmRN1mgVM5xTqJVZvyxJLsEler1yb2nOQ
PHjDV+4sZkCFcHXtn3OlOtBtJOJE9IXTywad8sr6RWrhFJvfNd+cGXOAO6WJ34BIgQoaqVO76N+d
WsyX0injhxVD1H8jGCttXP81eNvBDChJu6jhYBIiHIGIwqGU0Hbz57zLpn8kT/Ievq5SVxFFvhWW
icIOasCSwRNEbe+R5k3JAR2n4oYeNlvlXXO+3JcCQjvhSprEkZT4g1hQVX2nK83qKyx+nKvril+U
+xmezwiQRDxy2sbqooyXPIsjWIRM+AnUiooUmTR0+s1H77YPENWqMyJJzhBvl2tlzK3fs12T1Ywk
D3R1pWCLrPHwiatK0lfe9Yr7Vg/UVSPuxlEMVCO6vRu3FkYL/F71TZeNC9bpJOxmz68uwvtnglw2
G2lqQBzUEBaxZjHJk3DoASRYYj3R79Vid5QNWSIL3q4Asj3v5kS3ZrDucK/hYATJyyF9FmHNdwhe
spcfUGUxuEDAyklodns+wSGSUxLMgOdlw8NhCJWp5EN7oZQdVTANIuZe1bBgziSmN6l+dJIato+S
3bb2qWB3iz7LRqXc6Fg4IimPDFjBfmh8RBo4cvO4+qXG
`protect end_protected
