��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#��R�C(>�-|+����J;���5ǔ8#.5Ⱥ�`0���Ny,�iOK�պih�W���?$���!��p�n�d�v�O ��E��C��V͐+@�v#z��O-ћ)��[�����Du3k�2��,�A��#]�ɑ���N���C��q�$Ags�NJ
7�n",2�b�HI��u:�"u K�������� ��)��l��E����5�3��w^�w��%��%<��. f�˙�w#��zJ�=0�����@Y>��A2�3�V�&�6W�EU�y�
C�^}S�(B�h�x�g:���%/�(����J��>\�C�錄�_��gC���S�~H��������j �Ap/�����wR3� �j03���B��Z��΂K��(�ؑW�,�����\�^s7�x���I�>#���8ꦙ�Cr�/Ń}��<>>��fc�.���)�`�g֤Vt`RZ,�J{���
�x�V	^��R��� �R�P�W���v��(��*N������^+�1���!�@�6�{� �_4]>�Q�'�a��5��A$G47��kd
�ح��"��s�������Nu��S�n1�0}B��c6�����4�-A$S!N��ω�Bi�w�=�3�WT �ַ�2`����Z��[\q�Z�:;~��򵓲s T'�(@�$r	,��&C.���糗^m{d�mTH�n��CqiB(�W$�H/��9!�Ux����.75t8W~BM�![3n��8��3�[Μ��'.A&��ypȫ�Mw��FX�I��!���m���3N�������s˺cv6����G��a�A��.�=<��[�|�
2xT���j �:���{T�ґ��'ߜ1/1�Y��F�h����VK3����)�gD�UѰ��+���	���#����}rH3<�����3�hn��l��o9F��:+�� �O��k�nk��l�k��ŏcz�b[���{~�+�b�U�_Ldߗ�k�\06���T�I��LN�N@�� ׽u$�����;U�m�i��Eh��Em�C�El�n�0~�*_;#3��OuB�M���h�����
���AҬ����:m��-W�N�E��Tj4H'6e��*yW�-D�[�@AH�Ȫ)���W	��Id̸�p:/WH�>qx�w��[#�Q��іǏ�:*A������%�w/+C��O(�0$�O�>A�2���s�/�aR3ɼf���h��`x,G5'�b�+����e��x)9~Q��ɯ�����^F-��I��_���Mir��y�$~C>w�s�}�����������a�,�����@�;�<cQ��3{�����M��[��1�~�~toU�p\��i�z:╺#0=�q]�̎��7 E!j�����rL酚�ԸM�k�����y�<H~!,u�*1t�Mt�,��3-�P���:1�7�,?}��0��2E�����b�)�c����,� (���F�����Et�.�b7T^�����?4d��=����a��d�TG�M���V��-р�EZ C}v���6Y�c�%��mF�Cɳ{̛��%���;`����Ixo���i�_��LܟR�ܦ�Vm��q+���5Ѕ�DS����N�tgZ�:���-������ i����(���K���]~\�ې"�M]ׅ�@9T���Z]S��������O(�:6|[Kld�=~��
������#���4�|��<�~D��r���cO ��H���q��LS���� ��^K�{Y�(�42�X�P{�J�#���G���	�f
�b���U�fcq?�.�RǷ�!��^47���S��ϡ�YY�\۠;t���FT�������`��$���D��8���W�8�I&X�5��]:Z�|"�ZJI�>��H���xy�d0D��]�?<�`ba.���Y�U�����k:�C��͸��^W����T�v�A��h��LA/�>q!�P�;��q_*�,�<xX
�e'�g_v���'�"���j[F�&�p�OmI��=*!R!qŭZ�5��|: 5����k�߰k���ʇ<K3��֚�wR��o���[�ʪ���(!�if��4mY�F07j�����	(�k����F �yY��.UV�f���~�L�{��C���<N�$����F�y���;���S���0e�ד���1���9Rh�PG'kM�|��6-��LM4*���ia��C���z�J��`��1zg�&��<���;C|�Ca�H[��w8��w����M:���|Ň٣���SdO���������~�7����IߤH~��m���*��:}���j�X/�-hd5ڊ8g���b�B��cM��]���"Zú�p����}��+��^1�������Ir�q��!x��q?��v�����YC�(F,G\�Y9涳��R���u�EI��(a��p��/�6r�צ�P��Q`�l6�W�Y8XK�g��F@Ȳsm�<�!�@�v���^�>������V���4+h3����h�3��5�&u����#,�s�HզNSJ�>$��m�f�����$+���D�tP��m��\*_6��Y���z)#=����~�4⮶���=%�������M��W,<ْ�������}u�C*�GÅZ"6�}px��������"_��&`E?��}���!��T{�[p�}�9��d�72�S*�ye��d��s+���Q�^&~*3���ӴG�f��7�jL�Q�7�[ ��<n��p)
�(WZ����-�U�)�O���Γim�\v�4D�Rҳ��);úM�}r�5E�!��k�8R-�:�^�f��(�D���ӀZ�#��׈Q��ڮuE�:1��DT�i �[yYe��Q�%�9w8?*!�m:�8Ѝ%���`��Hd���UW�8
fI�ǲY��de(*��GB�R����`�'8�߁_���S��Ɵ��`�e+�&�-�����e���aC�����d��&/��qل��>�|����r�j3m8/�|G�mE�����h$Bº��%�xQ�y�XS��3�o�����'�A+D�ߜ�R�GL$�,P�}�@{@�ј����J��-�n����;Y��-�اiL��H��T_*R��\�e�ۆ����L�a���A�,F4S�-���,�	G�U}�  ��3����`���?h.��I�a�Mn����F��66]��߾%$�	;�r�m�V�kݿ3����#�
G�׼߬�¶w"�M~┦�5����Cnl�X0��m�}�N��V�������N�%�Z���(ō���
�� aA�,�7:���z�/b�lb;�����+SCו��ǫ
�2>Z5NuR�����GK�Uvg��6�1� _R�p�[��un+������p�^�r<:�-�Y���[�)<�+�.1L����ӑ�GƅU(�X��|�LWz�if�KJ��r�Y6_�1�0���m~�8����:%������<�����#o�r�͍e*r�d�#rVd���g�?lJE��	E���~"\c�J%%�;��w��tv������U.����a�G�4�*�R�{X�'�ݼ�8u�W%�@���.��Ǫv�%�͟'WbR��h�.a)���Β�b>�~���L��g6��-�bU�a�����;ОM�P�����"�9���.X�%�<��7���uv˨�hgurNf#���0V}�zC���0�#����/�oR�{)�մ2��uKx���D%'�e���MY�;t�i�3��$s<���&3��JO���sʘ�����D5�-������eZS9jC�k�q�m�O����4jc2�J�[����Oc˫j�ω���~�C^���h1܆ԅ���>H1����m4�G�� D�����/�Ii�T<`s��_�B�Z/��pK���mb;��� K'�%���5�k�r<)�,�ŧ����]�]�wȱg���:�X�~k_�{�Жo�+��xb)�	+ɠ�L��=�B	�z�5��t�/�Z5)8p�ՠsc�w�:62�w>bC0�|�v��FlV��5*�b*�%7�W�c���4�q��8�>g;W