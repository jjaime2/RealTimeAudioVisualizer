-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DawWpfu+4+XXWsrc/OMwIzBnV6FbaR+myMmc/HQxn2RGWJrSDv9vUiXEZmHJ5/g3DOaZ0s+Nxz2d
OSZIiHUyiWMtKFp7zAMLP9NnB67qoxuTBoDRNgA3no90tAm/oSj1HNMgoYltJTzCHj7XotE3i7m1
dvSByJr457LsH4cRKdJUuAv8Ulg6e/baVbHKBbCslbx0fRjKFl6LehMsXEjhbaDhmt/oRxfUJzI1
B9P/afRLh5o/et70XoRp/S0NPT+JlGAjnv+ZMgv1MrDAGE8cExrzBq9VVHc/hvBgAaPw82X/g+ch
VSS3k4PdJHxPSR8vrlXvx5C6r4dJ4nAKfy7tmg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7024)
`protect data_block
gvKSMceIhQ/T30g7PLdMmENxoeNsQ3BRczy2J3DjGzRVPcfCQfxyhE9+3G9UASZ2UQtVdTYo/1Bb
XBy+3pf4mzluidWpNCQTZsp7NZ/uKW9c2xCBEcG35pN/svUH/sMNUQqXx8n8a6AdGrp4jyb2hIB5
LLS/Ljbfz83JfU8Ywd5zXKC+MZBxzqCbZgVf3zibBlKTTMDRmsQabMu9jFTrVRhhNwePcINvVxFR
EGuNeLCqR4SoUU29MGPEqjd9TFllMHh82DqdfrFuJPnEftnfZ/ZlJfs85OMggsjTA+jrgGJtDBhm
mfXhtJI/o6EsKIdMNtLZ/xDyelUBXd68ED4IEsktxOZrkQAnsRW7zyOn3el1nlfqH3yZc2jd7By7
suuOtl8IALDYPwbXM2pXoUfyirur+f9oigfstsg5Gdu29/+vV+qEJVl0pquq95rjHyBEy0ZaLr9s
z3plpCC4wZrfpCSEtdDBT+RGLj4yPRXOqv25yQv8OGm/Am0A6OcpraYu68osPQ9HRN7/IQiHfNne
9As2T8Vat0aGM850zwnEZK+a2OkBUSpNUhLu7KYxxo3x3Kh4T5t0u6Jm6tVr1WDl2uYNsswdwXV+
pnaL0WyPCOo4Ga2ymRZ+IyiMrtSBk/mA3LXUjN5nr9CtYR8UqoUnXqvG2/zsWm8s+uLO9Rpq6Wfk
4V6OKUqManzN1nbwg4rl1gsKpVSuqADRTXeLd+qIle4fy+EngKRQUllCVX2SsnnoIWCGM4a9PODF
K9UfOCe07nU4pzw14WEisQVVtFKu1AxWJa3GqmA3oB3mGOGfJeanYbNpTlaDwE2gxR656kFNkd5e
HdEZzVMSjfwDAyNbf4ZQmkQ61Xem3dWNNzLnbe5bth32Y9YAinkHAT3MCI3nzRHI5bo34/vkddeo
HJiK4mfZbNjoGlrIEujy4mBT7NGYnfaR3xpEoMAdaxZuDekdN6HMpiTnvHCcy4LrEqhAxpIspSJl
KX22HTtv7gqwLYanF8m6IRB/u6c2LWBt4B+p9o/lcd1239IclaC5oLUWetYtgkxFmIU2IredTkms
tdyU6+Ezp9mtfLDrF0Ru2VtwHwxQjI1oovz4q7a/dmj+6EthTmzqpooCU9Zkzk9qVJQ6214fW6EF
MA8Gz7SmzPjKAW4vKIiTkS01reghGdtpS0onfP1nAbkdoYLw/i47dSzMj1MBLOVSOkhCNgHrQa6h
pI2EPEE9Bx4c5BtkG0BYun2oeCpeG6RumwUO/QVJxWU/lzlzYU3JZHOBLop2WICcDPpKlVLvRqyJ
LVaWZ1rMaLsZBObzdGQtU4BNxBGn+/Apge5zPQBpG0BuVgT1fbIlG5+kyirBaj6ZW1YpEvIDfm8n
2J6jChJefHigJ/YstHR8hAkccmswk/Disqsi69yJ4nrueJUwQdcV+pZPnNKQ04S5lFEJ6S8bVsp4
PiJpSQmCv9q/JeTmgNfG/TwLELpTq+43WWHh8VK4XdpK/eFYuLMM2vtlRdyY30Ze0oxU7ngNndLd
xDTqEhghI4NSO26Y94YtHB9kyU9x8Eh5cn91fpm0IHvbzvJlBF68w9bG7qc2GoC6pmmgSgFLG6CQ
nAufixUXpAG6cMP8Q1y541DtCAqpLFPlmWbE3W3MKRiI7XcJI5HmaWVwCwZDemk5YI8QP6OAKnUB
8g3gXoOmqBC19y9w4ijXzovnNQnovMm8sPyYi1+J7s0OfnXiSwAt0wPRcKVJUz1uUVkHYbKt38q0
2FbAceoUb1B+0xC4P+DshQ97r7H9Perveug0MPQA6pFuSMi6WcyXm+Ytm/79hpqu0MU4ntP05osi
W1Vu83/wUA0g3fmKBVgVCLVK9G8DEurVOo+pHqRra8q9LYjiMX43EC7+XL2xAqe65LQfUSAiB9k5
fDKVjjzB6z8ngGUQEqLb38fD9Fl+CgIP+fL7JnKNeoJbL910XNXFEmYEiRy1828qtFba2/Xbctd2
ljOIZHc3IR/oaNW8PnaM+X1NkmImDbGqj7Wyk+YPxnkgNqAiNiFXsGAYFRs067O5nVVddbZ17wlS
mnsXgCWDi/9fKJQf5p274SMYTKFV9wBzPP0jgDtcHUL3itYFaSt4FO09s1ECb1X/NQTGTI0VtaCq
8RmSI6y2zmmf+Pnn6c7bgczaf6v7OEUp/OFpcO/c5Akvj41YwEFHD9js+M8SpAMFKf9gzql63LtG
P1GOh6hiIAIG1sSF1vnpRbgJqhYEM7QBbdyUO+/9VaSdg/Vdd0iX8kM2P1OXt6NvErkTvPfDoU+D
NnVbmsVjs4G6MzKVEy1bh2x5lZVXTAeYEDp+tj0b4zwTlDOosbilZBv4KZSu8EW5q8qPSEgOM67f
yAc+DdQvjnSY8AIagaR3UEv3qXZGRrThcnoMsvw2YvvQxb3AnEHyVCdPueeyuVxxC5Gz2+1W51nK
lMia992cyt6+NPknNsthVAhxSoyCvVcAMYoCN9YJq1rm4yg1BTeNL1oyJ+94+xmQf4fxX5uffDoN
lIF7A1HM7ODB6SoHVik4lzj5+h6tvObqtmv1J0y9u62hSC/UtnFzgYeug7HOf5Xw30HVbR96OHKl
Kr+/vtkPnm5cy8D9qUMmOJWLzS+3Rv3ydaM8D65nBie/lKa+lrRtoJ03Xx52OMRsZ28ge/E4zp+4
gFZVKiFYio2ud0WcDR+GCxu8Ebkuwd5QifO6dkhVFct+YwOM4qLms5BbOyUhgxS80PU1XsfbAgAg
I5i6tZ1pIG6gnQfl4bIt2sjwAbNf4sEK81bLVNltg/NNkKUOboMfPWQ1qvdgeiOYzgqPXPv67Gz1
fulHOA5GViXZGnnkFTH8iaH8gYCsU1xoJVuQda5aFn0vV6RKpYY3DN7rCqQ6BvU39lnyINhKwWrj
ABU97cmbTH4KoBwdTFpeg2N5DBMp9tZR3TmJbBz6IJ0pTDkzoyC7YI0CMqYZCZjJXggplXdbQyNl
3BfN6dyjD16WIb3NpOVylo6VQz3NcTIQb+cxbEwvhhujXYk26DeWn6LejgoU6dIFpz6TiZLBOvtB
WzidinpGRL8T0eATfVa5Y1dxdkwzck4Z6OXdiP0CfeeNsO9gOfsgN0p1yVx5bAUTV6adPJu1FjvH
MA933bY7jYCh20TMj1YGePFubh2yYeTIr5SLu59RxHdUfQe2usContNx1zkT/2xasY1rJu1uXjwB
y5460C1M6Hj/CefnHBNzOsEWsEVxVaMaQMiLHu6IR0BX+4TPRTLLFwUkNMsPHO3rNE+U6IRz7tBW
QXPvbwDX35Yt2/lGjtdBYfRju8cZhNxos3BdFZbkEYI62cfvHpDSUdH7azaFuIHqHx6VczMEn1Qo
28H4Y8m3JZcNCjQBcIsEGNdbXcQAfp72oHq/0z447l2aTFZUdZxyrXyzHnsqqe+DeHqtkHxNu7Nr
tnt2wi8jZmAuM2UUOBYvIIAeh1wAfBZSk8FMoXIaHGvENwI837UhqmVFcqpgmTtV6wPVs0skZesl
FSIyLLWl46v+1ZmSWsY3wU+E6+LC/E2VmD9tvHDC9d/T48TqcKuAFsqaOCcC87Eul08mbhtYSAnF
BUwKONwNXppKsVPZ5vEPFhdGggXAh+fcFchC+Ciu5rDtepNAh5Ega4dYRtC0yOHoTSu2oB4NhmHD
L8gZuaEiQN6OFGe0sYY+q3JFsgV25iHMgH5JEXIvjQwqp9RSUxFgS6MdUCZeUJv0zP5ykodNR1Z1
VQ3sInmXg0Jc2JBSZdEZyeRhS4IdP7X+rYUxREYlfTT4d2iHgenG91zJR9RB6s6Va9WTsok8z+MG
ecjzRavBLSQ45bqbO5otM+Tzog2l+Hwk9qgTOVmMVZaqCZbQRlqYmDYEPViXVHLUDvpxgp9o3lSa
csTy4ovZxvM+xSw5ynH+xhFY7sN/uO75NSb0Atgon7c0N47Qehh/eo1phZ1RcHoRkv1oFcf+a6ly
fWOq2agxYBdWSiq6jlRFsQDyV7OwCkBEFOuQOYVc5bXCVfctAuc3yrBCIacx1co/IsmKaEh08SiZ
07UFrzIpCpi2ip0H0pGhFEF7OgVO0XaYQ7t/IOYo8tJUAN0Wy9sn3w9mMC0QrWywt7WJWZMMamrs
vt8QgeLmgEDThsOMGP/1QbeVPfgIUT09xHKz68C3gf0X+FZVNqYBYmawca+UkdV2yQraK6C5ppDN
8YLeNCv+8DC2WAjdiDiOyFJ8ifO1sxZ3S0m0iL2JFJfVXGX05LFah+rjCuBILPlH/kziRBAB5eEo
L4S2/cHvyp0Y9cqZQkl51C2stAOY4T0QQahu9ZhxJyi9DQraT0l3R6ZuREvrUaKVPco5879DkDKU
4Ub5osTvU6acz7qOHnktKS1aY18w0dTRP6hXj+is9265u89SP/RNDSWjqiH7khNDBIyZkQy2wsCy
I2fiQYBVDnt/LqfBI0+j4ibneIBppJtsZWW5RNEqD56OPPHUtVhL2u6cY04KAmqrZBSIWDy3o6zu
YiL4O848OptsITzvmz4KsQm/EsAB1VCkrLAB2jXSKjDB4NWwDkB138TVo034+C5xBNnUbNC0p1SD
nx1nwiOpn93qXy//NFks8TwrWzXFCBiNoyptXcRpvdPsJTbUDfcdAJIGld/PYboRmbOc/Ig0Lxwm
O2zzmWuaUe3XhNf4NQ0ZEQSeykQVzhBcN3563B8RWCdCTMUh0l+J4V8uFLMR+2iJ/TeFUzn8Nw3x
tBmaahOkCCIc1isYBhYM8w45kZMHYlCAH6+PaYSvovjZjLuiLcPjtVWLh6MTCTYa5Nclx3CuI31q
pYdJNAtmkCr+kjjE1TkDCFvAg83NUsQ0x9Dl2GuPMd+I++2xH7Mgoz1t4E/U7wWthFjVfSh/pKWg
e0EYVG0YS+WPVbC0MvnDbKHywNZG517gGOOYW7CFuZsfVYJx0TiYGsaHDDv1nXx0RUoqXYNcGpbJ
7ionRJFyJoeMQ+kAAsQls7x+ARR8duVfNEPg0lHOg9b0Nc11lcSQklVNaUxkKrHHpcURJK3N8NFV
DVtM2P49wgZLUFEju+uC50gyo5k5q42RyxsWnErKCB9+F6e9CgyJ5Jj2Wn4FSAN5/g730n2StFxP
aqVC1SLNsQOVnUij8bjf5A8L8YuMg5PueZC7RdHH9FjJijhLb4sKcjizItiZDhPReni73c5iVK6p
4Bp8G7en6StW4fpQmpHsQVYtiALsvaWNtk4ilxYAUPWXMY2et+8j80C3rsi/5aTaMT3Fs1hTbwHY
c9e2wVw73Au4Z7Ggo6t6eRxbA7jQL+qxOA1Bx7UtCOrnue3DVGemUgbrmXdQubCBqB+YCmMBx2PA
LQUkrAFOTUxhAel5zWBzVlwE/ZLa4JSvXZt9aPQwifvbH9y+C09r/llR4g29ty2S4tblfmtjx+/p
HTBXWRmq5eXPuHUSO33YFXebhSzAY6x5aGCi4atXgGqRtnJxrF7berxGP0f5jbr5B8c6rq4bIJei
GrazQFgrOV34WDLS5c/xXIq2UsPKnYOOk5qFNf+1qF3u/aU6h+fBO/olyWxQFapUcwf7jYtnDFFT
T2Pgf/UpTa1s4ImoO2AT/fV98xv4RFdbpUyhK9Wc9rw5jBOBnxQvc/VrrWWIiJore347vnrkMYcb
85o+M80iItOfFvUvUz4OEj9d2bHysw4x7z9qtuBjCPx9mqL03AAD++pJn/E1e4sothEVNb5ACPUi
qHfpYnKGp0x+3mDoHBdJ0DbJFjCEnpqEKHkmy8QSoVGPUUoemqqhTKf8RmKxDzY97NZdOXI3zR4/
OcUj7/avJo+eFFK4lof6vSqllkPAc0NhVGy7yyylnJ0nGrSTGFhxlAGyBpxwtoMxk7NtXRl15K/m
UG95yTwEDwr9UktOiqjPJnkfPDdlGxY6uNt4tfjtCWYi0O8uK1F/u8u72/u2DyKdBknq4k29epVY
2M/dwE7CEKAEM55v31xOU0l6IyHkyY9hDrdiJyjyJolVdjnQQ6CY7G0mz4PYsGGyoaYgP2Jbfwjx
tVrGGRaBWQ67HTBbSobbfpqRdXY4ihRo1JNcMowUvbyUnhuOBPNBdNd5abpsl+3C2nrgB9UH6+/j
NAtv6jzLQyhWWYVXEbAY5+WRjHp3iJr/7OhQylhzioG0smk+3scdLyxwl6cJNUnp7SBLyeQLlpLH
0G7bkeGunoh4pfoupGe4QYuL/kBrDAcWdePe4jg9e3fVkkolirtmEkViA+p5kc5R4MYahA4RtcBH
YhuQD4x/VUcI4VAbEdsnnS7ReXegayOmE2x8meXsYuM7PwB7YxfUKnSAaOMpMrp1bmRSy02sPDeq
29n3DI02FnGJojfOLo4qf/AUhCDrL+8fpdVrW7/6ELSdmZmMGnjgrNwP9eDeE3wtk6nUomjAvkuO
wdxcMirOaJa+dUWT+PfXXfLMw9tx3pBtvxGYOlwqx3vvoYOdhNd5WShy9GTDoEFXSJyZrpsm4WO2
fi8B34oEOGzMDtC/7aJCZfl5VJorpt6r5WB3AQzKk5BtvQ44fyQ9HZt3JNasIBGTcby6a9zFvb34
+jA0Z6ULq8D5Vvcr3XcR/8hJuNInFUSIeF/K8qgS2D9/d9xY3UC9h7fXHkbxwUwoD6KhAYC9Jidz
EZ/CNSFMQm+V36E5nXw0hHjhxOIDrSGv64aDl5taQwnYcXjuPCWnQUl7f93LP66OAxzF81HHrFgQ
71iWXMugtnh40u9vqC/sNI15uxKwhpv7/SDGRYo7gBqXF/iu2amf1sb0k7u4StQGySxFrIwdFPDp
9M/Ibd0FGysGpAAAs8cCKGXRRHIKXMJAeFFlqVtjG1VxfcahC391rWevkX7RnXkTnowaSHV+ez/W
o3s/ACCwOfqFBDF6G80hXCG4szHXF/F8FC7sVZQQg88nbASGrjaS8ng8hFPA1alTzB1/q5MSCfLf
bbhsxYsDg8CvWidBf4C2GzeNQDSME18TeRfJXvd1UcOQXrbPLLlLgkFShXfDYlOwL16CUU0OK3Bi
wKYBoVuXfnBAyyV4bv5oTWHQ4E84h5yJ5G68uGulSqgnEOgP6Xa5pT5iunVK3qW9eXCUyS1WSh9P
1b+WiCxjSuaavpqRB5EjLGTB7u3Xqc17FqeyOidW211jpWnJtBpL1KcS1GWl649a38cWZV7CXA2n
PD1hFTd+X2p0VdfBrXzSvwsZBgWOkuMJ4oxMkYY2B1Lnb5XW5gOwyVuwu1+uweTmo1F6V6dEzlLX
tBSKLSOAiwkO8u0XgWBv/31L2U4Y926Xwu7TRxvXBQ7AuZOQUDs18pAh1JQFb5ybJhrlaqg0i5xG
UV8Hq/uKigRV1zRdFRelz9Oqpa8l6IWMLkidR24X/4ktXFgDrdEGjE0Tua9Ry8xwdjyr1oD+El0J
7AFobcm4hg40GaVqWhoFko958pb4pOk2zdaGoBiFPSHTcRnHaCU6xe0NY8A5AhOIubz5vmO1bBUE
jBF4MM8qBp2UHdBaM6mk6OoR62bCs6yhiAkcmgI3TLSPGWx08ZcZAm4014kzG44FPRwa48pmsFZb
5vSalxpHOO8XepJffkzhJCNkBYYXv7mBXgJy6qxxqBdNheGXKDA64mtjAAVrfgvv3OSO8qAIUiSD
WMfxX1UMrruWZM7InS9kQZb5uBtSw06JC3/3/eW89q7ZbS2yIbU9MG8WUDLBJA9Gexv24aKapsUn
1YL1YUQkroKeeTr3gg8RDQvJssn941eJuykNaMaUUb1yGqaE88m6q1vVZxTnlOfHcoZg4sM2aGy0
qvf0hhg23TRQMM7aW4YDaslVfoCrVPhChBPCt6J5tV5WjVFeQMARPxpNnwwA9VpjvNfQ1VcGY5U3
DMp48Ta62eRneapmjD/pN6fBhb1lGeH7pmpKCZu/v06Fy/Kfd+kmALt36SGHwHUDX8lXQeb5JJCO
bQcg75KW988klrLJdV7hWmC7w4A1Kaymi5ghqmZGW5mk/tuuuC9f4UJjSuNw/ivMviijBF6Y4IPZ
MMaJZS8Oq2c5CS0nLf92BQ/7x0kWpoVB5y7Ol0ULDe2biHkC/fiGDReHjN/3lUsd4nBipI1GFgqT
HUWnlFnvdRuzLlCBMehUK/Sl73BFs/JfChiANmUAK4hVlSxCk1j33J7QC9syLR+HZ+L2mwJrn5tN
yE+PE/dE1XYY9QEyr3kSLZAxI5Hb4qex3Ps01q9ETtvBnnLAQNYN6sTsvXSDmFqJ04dvyAI1HvB1
mMiFKn3S1zaQXcsTYqiLVT3ssImsmyE9bCvQkYsd0d7ajDvPRk57/EJEQbMrrnFvtdCjlrcIp3+q
kxKGk8pkiYneUxR64A7WpXyhGgzZK+IbycqTnthoc25RHEFNRxKpRqsqAWSqOvM9bU3DeOUTHqvj
BL3MTYO8KYEkUmCo0EZ7LcKAsfjkSeN6p19clqURSxU2XqIM1ffy49Co3BPwMocVocy9DFD8jxek
OfIvwsH3tibNd2CRrL7e0WpTARXVqURWXHU9MnnIiAFthVH8tIZp3tHhS1sdeRIR3k+tjs3i2K16
p5eEWDR4hMHA1KjIxDyP8PKcQ1uLIwlv/+KLwnA32mAtUKt03AaGZtD6soXLCP6fRVwUyfwgB4Pm
8roirkUeyRAmjv10dOk8mhFErSt7pEc2Ias1oLb1N6WqUy2JxWhBp6kU+mtG93KBIl99R7TmwKS9
40TK49bQSfyr2Ps8oTADuAGMtCuPXtsiACvmwXYYEXl7qkqeqLc4sg644dyTJhYCKe64L2wl/UUq
r706Dl8e6Tnv+diZdqHsKCXJvKMVof1H9ap4/T4O9/jwtWgOqoK4zkg5y4JthbE5kBIhftiQYTSB
zlOfHCGUx0IVlIki+A/HTlJA+b3mUn2/+GsOzgOPuTh9H0ZqM9VZF/s0heLM68ObxT+FOEdqqsC5
s6hd1wnP0B1PbSrvMCJqbVlGB5731MEueJl7H9oYlCR4FTikrY5OrqV5ECtZsHICZekLsUppns3u
1t0V61ccVDywAwRRi5hQrjiFvpOXBmmlgdkfhP0VGi3MCubvPyTkcr8nGSPVwK2TUUy/jvEdsPpF
Dh5rTFrrDgzVfJRBx8FY4oUZB99IxNYi4bdwF2uADaMMWVChdJ9BoaefFq1n8KHcJ9wZsdPmTI9C
lZyrmRckbJQEPc8KySIBKpxKq4VEGHQWqqZvpIVV3TPGouY2UX7wj1w/RGEtIFQhZbyolqaS5LNg
e1uRyEOnvEOaV9yIFl/r56xfkwRqOUqTqtKwVfJVR8gOCddts8Np1Ec+nriQ01L68744ezyfSiGR
zbp5BMEgOSIn9ERFNwlLUyeVIhyFV9d0+jArKkylQVcAauOl92E4++A3PTRyWjM2UozvSLyl0RZv
LJ//oJY4FyPICQ8ZYA==
`protect end_protected
