��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ��(w����E��}�U.��K0��m�A�x�����m]�ǟ�������"m81T�A�q��z���7��M����~�`�]����9�Q��qۘ�C��
�'�//T!�ѾbA���sq�]��[����A9���:��+�<��s�A<����?����C��A�5��i�NV�V}�������X�R�R�=���\H�2ŝ�`tw��	��v4(BT�����:F�Sݼ%�+�=�1a�M���ދZ��q�7�/K���:	��&�_�V�V!.6?(S��o=��m�4��X3ϥ	�6��ĸ�����&����2h�� �la�|U������F����s^�?�\�]2��8kA���lX�6�yAY髧�lL����vDEip��:U�6���P��ci�fPäz_x��=e:�1t7j������Ƥ��z/���A�@�:��u��V�ͅ�a�r��ʚC���b��J�[�z�d&qi}>������ �4K�]�ǯe��d<M(՟y/&�����=���M�����s(��� �F��$m���eg�9A�Oӓs�1�0=%�[$;�tu(����-���-3!>dx[�A����	ɼY�lI�߂w�:>���f����s�N�N����گ�d���|����d���..��'�$���E0��⛣��v���fCDΖ�~�imv��-�l�Uߥ��>�p�mV� �7"���x4抧���P�}>0�s�I��;wo��S����r�{���4������N]�@3X����ʵdzS2�4��y�3�&P��L܁6���M�	�OA��1|������l���v��t��Z�pr���tQk��h�,�b$@\s[���K��̛]�=�?���K�=|�vʴ/6��$)����&�X�@�fe�gы�3���nџ)a8�ͦ����kVe.x:�ƹ]bo��镬�����&�O5s��Կ����d
u�Ɗ@I���D�ps�,��3G��p8���#m��P ��im��
m��ft�R��`�ܚ��G+A��B�����h���8��>�D�`�]h�Yqd�B�`��0^}<���J�$���&���/����!j���� ����Ɉ�D�낿���Y���eu?���>ă��fmD��� V����8���ڔS|I��1�Y8%c.�m.G[b���9�L;��9$����^%��K�*��؞۫���h���S3�1��ԍY��A�5N�t��=:�/��I��|�OE8�Ic�|���:8�+(����\Q&\�8`0rzG�zf��[-(t�{�kZ��[{/�m�`$=�8�,ٿ�%��p��Қf ��9f�3yY�.��p���L����:��-�C)����;A�j��4~��5y��]��Y�pOq�䚡-�t��2�~w�KS�5 �u.I9�=<�����i�wv|u�dH�MI�����҃/oG�}�"� SQ�z����B�P5��Sj^��F>���*V
+$��^�Q{wSKI��n��-�l̔���Fx@>����;�a�&\	�����<�Cjm�|sx~��z0Ͱ���S����(�쫗Gh0NN]����W\���ݧe�L=L0�m�LR������>A��̅�{��{<�[X�lc���0��}(�]p��D"d�L��i7in��yE'X��!�Y��	OO �9���~OՏ�	Ѫ��n�Զ���W��pyކ�)��vr���?��zƳ�I_��D��,�����׊�pL*Rj�X�̤�:5�LWTY���]=?f�}f�|�PfZ��:sY�-�m�DB����z�<�Wt��j��[J�-��{B��Ӥ�S1�na�������U�~�����0��Sh�b1bgr�ă3�"��eܞq�"xsقv��A��e<ȿ�_A�o ��v��q<W_�������C����wM�wI;#@��s�ёK��P�Y��^���F�C�D��ȥa��I��U]��y8�6�w�v������7��M���	��|jOZ�u�;�����?\���jX�I���W�4���3.W$9+q�����\�VoOJ�G��a�K���@�`e��ed| ���s�����+�ta��.S���������k[��Ƚޡ����sk�w�r�cͿm�o��
r8�����2�(��W�Z��	��{���tqmNW��O�<��Y�V���N�����~�`{�\���˱��$�燹G����B��?��s�'�k?#0���L�QX@�T�T�������ێl���������[�9;��cA��7Y�=��]�k�yS���h#܊��a�q�}���~i&Et��5tL]ˎ+�Ǿ}T݃��Gh�&�/��/���vP�d���F\a26������ ��>Ԩϝ�v����bF:��������>��8o�� B0�+|��PPr�㴅3g��$D,܄E;�bʆ�g�%���A����iv�~8�|4;����C	�ϟ�[�*�:`����N��1�``�zFSԚ������7M?qfn���i�Z��1V���ez2�X�CX�M^i�bnGӪ��CuK�RP+d��*:�\Ԫ�#B7>cM2AH�Ҁ�A�15���8�m󆦨����<f���m,!�`��]6h ,8�����(h��>M&O@��~�:�g��2�6�)�.n~A��ԃ�P�>D1g��D��L_,d���5'�q�q׼p$MIƑ�	��l���dw0ZPW��M�i\ʶ)P@�+a�Sq����-D���y�cn��n��j�����Dc5Y��s����Ԫd���o���H�[�5q�v��]!�a%CS"�a�J��x�')a�D�p��>��2h�C�}��:�x��
�5~h�A����J��.�_�?펁���tc-\�����5�4��uK����LGP��r##Ӥ`H�o$�l(K�+&P�B7d��i�c\��MIG�5�ޮP�?���)
 ��/�+S͜�Y�Ќ���g�p@q��')�.����W���r3l=Ek}&J�+����A��N�������'MIeX�i'��,^k���cD��|o�E�Yy!J�كAVJb#�6nŇ��j7erd��R�:q�]]�Q�j�8��xh�VɁs�)��d�On�jr/�~��)�e&W��4~8���H�٠��a^���x���jD�r���0���AHy��v|���aH�m�%�88KUآs�+vf�(m��ϛ��u�����F�;���Y0v�W�1Q�h�i륟&>�ʓ�.#�a��뙀���$Gg�'-g-���b���&�ڱ>�q���P�88h�n|j|���z��E��?e����uY꧉y#M�Ν�(&t�+�>vI~�&TL ��7f��쵦,Y�x�J��p
s���Z2�Vh�� u����+H���XZ�u�3������nժ3�R���$~I?�A���9�
	e�v����H�9����W-w<�x�G-&�sE�nF�b&��S�*����v0 �����`��ٷ���u�|f��~�鱀�=�(��=V�~���T����=�?=�^���U��7��>q��NGYFY��^�M��$�̲ZD�b�M�8�wxC�u;ݝ�1|8(aYg�n4�F�6��]p���C�"B�V�P�)�."z �tc��q�Vne�8M3\���P����HA8��I�J�P�����l��l��r�j�-�m�� M�]+��-*�1�����xƞ �z ViK�_�4�;e7�hoQp4ػ^'�h]��.���̭�92~�!V	Q6a�������h���s�j���_7-q�����x�� �}�<b�� ����vP~�S'����j�ͪ��0�6J�Ƶ�t��\J�b��h�xk\���щ�( "+���/w�q�`��2i���bP��?�G����9OUM���e�2�i���=�4}f�¨ԍ�e쭜#"&�؃��� p���1tZ_�5�kfݩ���h}�RcUG�вf@���B�������Q�N�wwg�n��[B��Шڬ��e�'F��!�E����R������J~����5ꏼ���]�D�ȥ�\إ��-�8�snѯ�m	�[/w&��R�@LI612hﺈ�� ��!��8�D�HQ���ܾ�+��W]|�����v�Ԭb�6(��°���'���c2��g���(���:���/�<�O���UE4��w�>٬�v�9����Xp��ug�lf4-���d-a�daY��9�e$�[)�p�����l)�p�R{ͻ��-��6m[%G?�v�o�vy �.��ln� �:,'�]���q�Gb@&?x6�q|�����-܄�s��|E�fw|i��*��<Ú\ kNc�a��y��YU�i79RY�wF)�F�X}���ysa����;Sp����ƨ�U��EM{���%���cn!��n��G�$'��.s��>ܕ�A箨'�05���9HPT�u7�XOc��;�ƙUn`�dF0L����g�bؿ�1�?:����6֧=��7 P����P���a~���ҢD�\�~!L���㎖8����{q��g�ϟ 
~w�������fD��/G����+	�0݆�B�{|�յˑ$��rif��=��hsO^�m��&U����"B���>��_�ӛ��Q�M^G��5�~6a�Y>�S1r{/�0���n��}�}��0E�#�xB�)#_N0y����lkY�t�T�?-o�=K��҆�Z�w>�SB8�v�n
�B��Kr����#�9Y����?�RwuGsݯ;?�UI"�'F!�̑ɲ�x;<BM�ï�W Ѵ�1DRK�X)�P���<��p������Uf�W�0� TIlx0�W�,�g��-%�=k�ڽd�:�	����N�#ݠ����Y�J�_r��I���˒��Z����J�E(%tĸ����*�+�C?����͹�U��'��łB�3z.��q�7G*Eݖ�=�����g7���y�P�������MZ��b����&W����,ZĿQհhEX��9և"ӚE�vsn객���6nP%<VLB�bb�t>�c�tܣ��T�bay��.���\�Ps�|�!ݭ�:J�o�[w����3�q~۵;b�m).����)����ޟ�{_�`c4�����,�N-���6I��{�O2&]"׆�A=%4Hd�%�$Y����GأT���Ѱ��7Z/�IXt�&,�oء��g]���*	�-� �^�lw���bT5��xW!��k���a�Xҵ����.'�J&��ZFn�u|GK�`+��#��D��-	!'C�-i��l��ow���}OI"���,�ì��(�9�X��A;�CM	m��������}?��p2����̱�E�׸��q��~^�T�N�n�|�-�R�"b����(��>G�\,��[�d�ʍ%���+t���wP�������T�_�Ud�ζ�KRξӴ��d@��J75���r�;R�`���W�	���8�L7�	�,d$<��6�N>�fj����EfTm$`���U˛���]�3[F�QOdI�Q��������"Z7�� W����E��'nS��,�]��4��˼H�K:��]x��KT�v�i��~u�1��Ua��֋�M�w
��ra�@3¢*��D������9b�׃�\ʎ8�GI_Pv'�A+7�%����ϔz�8&����6Ğy�~��7����τ� ��G��[���}1y(=<���E��T?Zآ�T��G�ƆY�0���}���W6T`�~���l���D1��~��	�|����D�K���X�d	�e7[b�=twG�븺?v8�GXY��J�Z�Rn��Ho;nlmR�,�BO�3"-��C���rR#�oyd�`�����,�Q���R�p��ʹ�'��W�pt].�R[w�z��h� ��[+���@f*���.\�����G�>�(�#-���Ae�^�<�g�-:�ޚ��қz����,�y�0�Lp��' �D������֊<6���	��4#��n�bM�5�tlLU���&�#��y�K<aۦ���bƁ�ܝY� �,�W���@1&3��O��B��ڴ�R20*�'���ui2������a|��osm[�.�W&�y���ChE$����'+nV��s�a���B���]
Ƨ��� d�g1}��Ć��ћ���clEan/���ܪ�v��@���xA�=0����3�#ʥU^���)�]��b<��*�������=9"�?���0�v<�h�w��e�$�Z+R����V�a��Ț������~E̚vS>U��ͤ�'���$d8���s!����-�r�]%�Md���Lbp.�N�$���3��G*�Yq��1F.�Hє��3��;d�uP/����<�u��hP��J����QD�V6�
ۄ���MZv1	HC4bż�ﺹZ�\JCGB��	4��fw�+8�-���
�+s���,6��oh^+�ˍFb-o�>���H�<���㟗���G�AR@8B������e�>p�w���xE�@et�<Le��s6Y5PI�~�[-q�P}��V�̤Ok�~c.�JV��&�-�d~Ԥ��Zr�R�\2�g�.�u���-���]z%V|����MΊ��m�3��Ş{�Nȼ�&��Ǒ��,pd����K����¨�I�]dLmP�y[̄8��4G���׭�~���e�ř��a(e��x�}�{ps�EK�x;r'�^��ٟ�&�4� wA;��� �LRB��ІI�
�����&"5��G)�a����3WS	&�7D�_fV)ڷ�O�M�U�!@�\�}�����p�������`��ނ�#�3)��u�t[=V�p��q8&�Ro�r���u9�ɲZp�D�_���VO�b �T��9[�ana� ��S��)44p��i���3X��Y��� ��ވU�6<t��Ŋ�Ksz��ڭ�����ԇ޻��z��-+���x�X\[��ɷ�q�]p&B���ɗ_�����Z�_G
�>��<�>�g�(�������70��q�<m��;�{q���h9lv��Ug���Y9/��@��7��Z?�L˞7�7х�bva�V[����ڑ0㞴,LcnK!Sj-��R���?=� ��龸��CJ]TLԞzN1��v���<��i%a=l��j>�,��w��m��W����Ib�[b,e���H��r}�N�"Ŏ���KK>�f��p�����7��8D1���1���\}&p�o�%�}���U��~il�����C.�z�`�@�DG��6�vBb�wb��߇}�c2�
=:}r��ɭwmcL���b7tA�,�kg�8R|������!T�<t[8�v��a�n ��s����ɔ�$���|���<�a�\���)3pT'�j�͢p�<$���U�_�{����=���<F|(�U��(���Ͽ� �����V���9�&��B���!?4d����5�}r�3��v�5�Sj$��	��.���&��te��p��=�?9Ú�t�)Ya}Z������Ē���������_ѫ��؏t�=;݄s�aG��vU�}�;��'� ��gݰ<�V"X�����m�k�2�<&SeH�S�1��(=�p3H)e���������=���S1�T���57\����zs�9�fQ-DZ(.n���������q�7��G��S�	NN).l�� ��˰���*2�w;*A�}
�X��n�N�s���������pm��)n�#�V�]	���uያ�,�u^ث�@N����M��ǃb=K��v�w��>�1
�+.,�	}K���(!���Ɩ]KI|�9��y[�2�u�=kHr�{CM��3�|g�+�4#im��ͯѧ7�W%�N�*.����a*�\��ۧM��G,���~�f�+�	}-���&rB��˪�������m�&��d9�h�DC3�7�(�X\s|��3����蔩�{��e�I坡�W���������.��?���\�V�[�!�Ͽ���owl�Vjg>W�Kԍ+���(��rB~�XNv�ж,M�tfŹ�q�$xL"���������)�e���7��n:��3��Ƿ)k�.݆E��0�$��$�uP�����5��������z�ɻ����q3�9��F��G��r������49ݺ����~YϭᆣQA=�G��BJ)�^t�aA��Hco�r���(����n������_�W�Eր�I
m���>��G���*�e>6�iǊDJe[��	B �m�QK��2��T��(���at�Bgͤ_��@1��asE�}��>�������m�&�b!���y�4�~F��?䀱��(��I6���Nf�P���T� )�����&�O������Us/�py��3��l�т5�� ~my$u���U=��]�م�X�����T��M?�L=�k�R@?��6�1��A�<J
�w "jtZ�O?��o_�@~���[��|oP�s�h����FbG]7��)(h��=������Xj\�)G�Ӟ%3�i�r4I7����'[�x5t.�m�C/C�s�>0Twl�(~C���oGL���Ϊ1�>Z)�;�k�8�h�E��5/�~���� �w
�= ���#�����qU`&v2ںO��"e�t%m*ތ��(�������׃1vl�0�T�Ӵ�sSJ���kP�L�zB����gp|��3!h��]S!��[+_T��g]�
�z�Rt~�kS�ߍ����i�C%A�� #�2��>��X�ïj�)�aFj9�����>R�i�V�8&l��ʁL��S���-��ϡ��yH�j�
~���60�r?創W�TK^)>�JM�;�3�Ѫ�o�z�F�Ff��l�m|�\/�����V��w�@
J>���*o���z���:\��M�n�)YU��	W�[��O��-g'�&'ZH\�����jg���n'r"�on�����N��?U��Y�-�)ɬuWL�xt�PF%3�	���:"�"$��Ȣl59�T]A,fcBj�¦�t�����]��&I��ꌇ��?ϼ����u�L��;����D�[�<�X��2�R���Թw�"cQ�yV���+P�Ѧ��-k2�*�%�8Z0�.:����u����#G������C���o[o���K�'k��x�a|��u�JB�P��.k�����	W!d�\�ȩ*�d�+b;���a��M���)�q��eʖ�IAF-�%W��Nޔ�#<p}�'8T����V�i��:!f������� <y�Q.��4B�e��n1��v&
���Q�l��'�JЊ.�y껖z�s?vH�>I�w��9��>\����R����1��ac�ȡ��Vk�\�w�f�ϡ��h&-�7��;��s��d��w��ׅ���δל���5�x��ӫ���,�q��̯jf�U(���5�<s�ޜ�1�-E�R�?�t&�$�*%���0 �o���9H?��nt$�0\�6>(ū�:��"�N{����:j���E]yz�i0W򳕤s���9�(�gS�\��)A������,J0V9������s�?������1T1'��@e����}��t�}(��]b/�[�6�2�:_��H�W�m�S|� C(�M�D��$S	��8h�Lj��j��s����H��Akva��k�w�^���0}��}?�4�6յ� ��9d3�<�T�酜X'�T�b�ҴڣTHB����#~κڧL&5.-?��L{��z�>�3��6e��o�B��������$Y`f]}R���t�*d�|����J	uj{=�03��#�����=�>�^C`a��M�e>�P`Twz[�6�pe%AdEc�T��[�M*y ���!	ơa���:�G믍���ᕜi4��
��׆`���%�g�[坋��?8��KR2̽6d��˺�߅I���yn�b��he����5�nJr}`'"���U����	̊�b)��-����@��D;/sg2y�r��C'��s�o|ꑚLԁn�)#C�p�k�ʳ`�߁�z	�ph���/4�&pgA'f�Ԕ����sp�0��}пo4Q���8xx]��*�@Z�~˪������d�l��.G�6�t��g�nk׽f��,G�?$�}.�7��]ɾ$&�}�#?{X��Ɉ��	J��1��T`,�SO�*�%�ܞz�CdkHݕk+ �Q����SH�{?-�֘�!�������MBzE���3s~��?��Ȯ�f�aͧ�=�ꗞ&��ί*A��_���i��~���<���k��P]�vEb��2�Â�c3Np���t�t2���� �`�K7)��X
��~���*�@]ʙ:o�&�Il��o���1�8��7�T���I��5�x�Uk��?Ϻ`���`�ؐ/P�$j���� �Gv���ȱ��SUW5�K&��]��UD�O���������4��iv4E6������5ܝ�#P���\�K<N�t "�3pf�a�R�[@+8�dc0��,o���h8��͖ɗ�Ѧz�o�'�����3����lɏ�N�5K�]H������dj�v���"�I���O=�����kxǁ a�($t���*.������6ŌO������lɎ�q��jc9�C��O�&�[��|ql���{�ȡ������`�>�T��幍�ߍe�=3U�	�*$K)���Z:��RM�r7}�6͞��2&T׊(���z�^�f�Ў�@N?�7�����k���(���S�1����.f_���"Ɣ��q���h%�n���9�SB�#ź�����C���>�����{�����t)Q��ω���`q�[}$�ͱ[��u��t� �lԚD�O܊���noۢr6S��X���}.�\M^�.�F[w��NѮ>m���]^(���<@F)����,�,gG�2B�Q�-��*� ��쐆VU�ժ��&#{�M�Ā�S��x6��L�Hh����"!�l�Jk�"�01�1�RHz�r�:�����:8DthB���=������Z�@��5���,:e��*�ՅI	���_����s�*MUS�krp��B	�Bs���n�#��Q@.+3p�_`A+��Ү�!���g�\S� X�M���U�����-Z3����#c2S6��O ޔ!�:Ѷ�.b]3�е�iT���!��u�^Q!�ߛ3Ilt�A��Gj�FŹi������O�Y#�v&���Ŕ�fkn)���7V��8��+��,/�x���N�j
�����bҿ���w��x�?�K>]"�#kqQ�fL��I&��faf��pP��;G�s/�+G��F�f������gހo ���n����g�6'Y��"A�"��q!���r}}D-s�=�����J��(��H�����3RQ_��~w��0.8A)Q��aLi	�<�K�$m�W�u2�-�H���U�e`�dj�6B��13�bB/����+F������?����K�_��v�R�[ݳ �73q������n�{'×��*l�|$tٝfW҇���c�F�$����/��aV�����4"ͧͥ(|ES�!�z�#�qa;���m��������]�[K^�u��ct݃D�3 rZ�"�h�4������a:�}:� ����8T���䬢�tF+z�y���Vm[�=��N��n���g$��	��!6di��޿�Q2Ə\��jϓ�Uw���3`h���"��!�a^�K@�q���H�bu��E�:y��*cT�rw�����4�O����Ïz�9�e(�uJ�����j�p���x���,��N:*>�n���d�9:5UP������#P�̊a��}���^f�(�j_ᝩ ��ߺ
���T� �3�ݻd2��c�7o�A9:����a��^}*���ZǶ�,k�7��%������zZ<w��E�z�����G럈6j��� z	��n�t[�ۗ��*%�g"��Rw�ND����I�_*4!����0{U��(�:2_��y�A��B
�G��w��\��=;��[�Cw�C��ߥT��.��|�4QSk�$ή�#���L��C�"n.P�G��Z�i�+��E>�G��TCHT�_L�4�ܲ��[:6|���W{�S ��aF0_K�q�����KV�Fn���ܤ�i%�v��%��G�Zz�:�x���%�Ey��k�a�kqFKJN�H���2-p�f�!S:�r�Ĉ:G�w����ż���ῑ�����a���
	cȆ��ct��;�r����b!�@��KÞ
�jKZ[�y�-�	ǚe)�F�K"�+J������zh��|��栰�Ē�0r��Q̓��=�n�z
��Fbl=y�->_��V��=�X��ޛ���Y���%}�w
i=�n�Ԍ�/K=R`}Ówܠ[�O����#�K:S<	p�R�-�Fc�I�5�0�^\j�8��~h.?����R�̈́�#4�8Y���ʐ����ˇܺ�Z��9�0��+{��@�mm�؈
��H>)k�l�������f�>I�����&y,>b�+IS2�qmjh�ϬI��h�!���O�'x��$Z4��.�_t���J���0�ަv�M��3=��&���By��Q*SՌ���ott%�=�
c쥆Ux�U�q�(��/}���UF�I��D��EUSӓV���&tu��^�^�2L�4ֽ������JA�bv Tj`h]���z��d�β���m�W����{~u�t��9�@�����`F8_W��֚����/�U&������Z0�ci"��C�i�_<�~@��:����Б���զ

h�C�\x㝐Y˸Ɔ�+��HA���g&k$�8���+�N�(�&4��Z�"�z-�m�-wyzxc�c��*{3�8�u)fIΤ%�%�q8�(�N�z���-�H��Y�<29V�`jƣs����}ƕ�V��ۜ�b�F_�hM Ç4��i�)ua���NmY��@�ů��-Q?��%�n�	�v|��`�����^\SԊp@m���L	?��;��M|��E���NA����.��	E�y������[?}��`���y�W'a�A�00&���.�1��Z7���Ly�-=��]�С�ʓ}ÎM�1��I�u:��u�x�9o����{�JQ�����km��i�s��@/eۯqT����=6U3��,�a���l�S�=�K�JR0�+O���#�d�GE�w{K�E�S�|��}#&���Pw���lg��qB;���6W}�7J�����gT[�N��R�L��1a��
O���c�=C���VCDsd��þj7��MK���\�]8����e��|�nq!��;Ő`��0�ؠs��r*�o���) �#�n'��St�W���c���I����J/<G5΍�1�&疅bu��b���+�Ý�C��������HV
q��aX�<���)��gh:XM�ys4��e�n��f�=�%��T	�;�bnc+ee�*��A�{��,���S���u�)�~R"�Q I������h|��ٌ��!:�C����n��V)[���s�,;Sm��C �f�8�^yc�s���q��w��2�`/�v����@қ��a:�=p+ ��a��O���$�tU���.�����cn˻���v��^�
����L�L�#�5HE����htg�'�gQ�)_�Cdq�B�����ݧ�K�6���)���✲���!��ʫe�{[�<�)��D��7�56�`�L���ַ,%y�+���po���lҿY��v�N���9��)�Hg|
J�WTR��X�&�^+7y��wb���ء�%Ҕp���h�p��t�4H�G((IB�l�KG��S�¶�,v��w�	3Ͻ�����2H	䆋�R���ŧx��|���+�ٴG���lPiQ�{AɊ�ú&MD؆\|Ju�W?ߑ^5�^G�7���bQ�%9�����'J�G:q��>Ŝ���V���l����������l�t"��c_���P����Nv^�K�����;:bPԼm�V��x��V$q�p�����+������-��lR�ŊePR���.���g:h���v�(�v~S-��,�y�ý��bݶ�E2��&RS��F�����U?$�X#������0�������G�_X�)X̋��Au"������)8�� �����?m�^2e�[B'���፤][���b���	�z���p�z�:@K���x3aLj��|/��f9D� qQ������5�YS�u��/������yD!�ȣ�3����6���.΅6���̺{k��o�CI4��.?�>��3�7��B��ߞ,�\�f2'��VZ�;#�����(���!��,�d�@�y�=�g4>l�эm�Q2�p8�p�J�V�"9H�]�����U� c_�>�P�:=yv����j�g�r�ƖU��h�s��G.d0�9�-ѓ�[J��t䛁}�f�w(`x�qJ]��%���4������m�e��V ��\Ќ؁$#���ߤX�%1b��!���ce�L�k�_k�٪M:�8��`��z:��T5 �3�aݔg�j�"���w�وmm h2x3��(��ɔ����.6���^�*=�Rw�Q�����-
K����;���HVa��o��	ZڷF30Q��x����S��r����¨p�C�y�jb�43�§�߮m�zڬ��b��S�������KA��x�؍RU��e��\qM��+Da��J��P�w��TGmf�3g;�19���;�$e�;�}=�4I�6�(�_���ƕ�%���!�"Q���FQ�"u���\dHgQ$���8�AB/�'xsf�E����D�Oi��k������=�4[�镪�4C� ���  �e�`����[4j�E2T~�h
����C���3�ٳw���fW~?��O�kQ~J�C���k/@�U����+��vIW�CO�-V�Qԛ��޻�A�G2�x�����j����v���͋��ת�)��z:�`7#ꖩ;�� c�@GI+���ٖ*����]�MG�7}��.em~�ˍ9A�TA��|js����ۛL20Y��n�*G<�B6=V@1g5����ʁ˒n�IN�m����aA���qI�w���9n�dY�f	�I��G���%8�#h�JP��T�Q�:ts�I-n5o5^��\"�9ϏF�m�pM�e9#*9f&�fġ���<�^a� �j�����ZQ�
��F;6p�g?�8Q��T/�m�����\֐�yi���b�x�2l������\�O���.UQ��.�g��;���j5cO��t-LL��*�ɫ���H(,�1<J�Z���禆"k-�}�V�oQ[,l��`J7�Bp| ��/D;��k����P�*��J�g+�9�5���ew}2�*ؚ�ש]]jA�f,;X��o�&���v9C�^h�l����(l+�sIY� @P;6���Q@��a��U�j%:���P����Z闇�K�2 ��W�M�ϕj�������'A��]M@����a���	D�#;S�fHD��)���	W�[�D����4�Y���J8΅Y�pN�dD�{��'��=���^B0y�PG��E�+���в�(��l�~H�H"~�7M٧��#�7���q����S	�p��:i��0֞���b�$���d��`7x����*2�;@�����y�+�풟�I�����o�> r�^m�۱:��63cZM�Y0=י�N�V��r�$�"6� ��s~���^�	������`�VK!��Q/c�tp[�sK���w����*�CDz��i���/lnQ욡q.0U)���ƾ;^�Ҝi��Od�M�+��}�sd�	�����P?��ƳE[�Tj8��~���������.4���o��1�}��8�j��O�1����%��L�y�&  y��Gl��K;��B�� Y4�� ��:�YL�C�q� �z����w�D�>��|�i���i���Y�H���������.���QnBS{.^�X�JĤ1��4x���y�xuZgW��a��T���Q����BބʱF���� h��� �0Z%�v�H�!�^ĥ@ୈ�� .R�r}a6����O|���6Wj� c�Y�Blsp� ���&/U#It>��Ϊޞ�T��}i�8�ݠ��Ө9y����A*IaI4<v"��r�re�~d����1���qpt��w{�k���A�;y7x�ݱ۞�
��s�Ny#z��#��gI����[����Q�M�/�Y�UM���e�{��< ����
&�'��.?$u�7��2��Z�$�w����%����ě�W ��/$J�+]�]Dt_�eծ]ȎŶ�5|CǕx.�%�V��=�W���[3Ԩ�m)9�Z�K��.%��������WWd����M�_Fw(���BZ�+g>�!�6���拨.���	e3��o���"����7ooOi-�L�N��H�>���%�mo�ѵԵ�{�cu�T��w���ؾ/C�;�
�bm7X��5�������G��
h�:^ch�'�$��7C�t䱡�M��>���a��B(��wa�ܨ:��GIɱiN��a;}u�e5�<9�h��V���:���P���9T]�{G�K�º�I�~�5�>��c���l��E�("ar]��Z�ÌW}P ��H�j?�98�`%�_�jM��BD�X t�d�ٝ��e]�;���I�b(�H�0��o��L(���
iXUK�����U��L�`��W�g�'bC����EAY�WL	�nEγ��Q��ޮ��N��y�0[ 0x�W���9�^���4c������/h��0p���"^�V���#�b3���[���8�|����R�*���uRc�}�BSPR��w���a���d�����5�����߯����l���G��hN<H��6���Nf$E	�#.��Y+a�&����H`m(vk�qƺS;1�d9�!h�	��bH�fG���hdEgNG
i�!���G�`&�о�$P��nF`�ӓ���{�=�#?�������
�_��<BGm��O���~����^1�b4�ԏ�Ii�肣��!i�8���,M�5U��I����f"�Ca���k�ܘt�J�Wu�g��D�פM��'}]ۏ갵:٬@SE�ط%DF��rC8����Fрh8`����c0��s��Ew<e:�^e�����ךzl�Nȳ!��r9's����-�T���Q�H�]o�Xr�@l��f�� ���U2Vv��z�	��?��������J�����MĹC�S��pu��������wٗ�c��=�5�[�>�h��2��g�k�>%|�����i��,�B�b�Sд�Y�aX��)�٬A�?kXք���C���8����w��������7M�!�E�~���ڮ��yV$o��]qt]0wG���ت����P��#��I�(�|��Vo�2@2���u4J�NY4�A�mY@χ�ߺ{���O����\o!q[,�er�M��>Ϛ�Y ����ghlL�������/�����޲���Тmg�e�3J���ҕ�(���#OSP���/��?���UbT~���}C�7n2�h/g��qx0�r�,�l��eΚ6WJb�|h�Cԛ;�a��-���d(�W�l.��~�[����t�jc7%:��9d��(��$'�0�ʹ2�� x�ъ8ُ$嶐���Tof�P�[��hL�0V��9ԉ�euT�m��@b |��&�� �V��.8lۏ�v}�$��J�f�}SUn8Py쾸;���D�UM���y��P�P�l��M4�C��е�"rx$���=!�uԶ�� �#*��Rt��p�={.���Of��"1v���v�*| �M����K�r�۰,��UcLIp�/X��ʘ}���%Ҥ�d̨�0�듉�3��P��s�KS�j�[z��bG}��i𢾱��hJe<~!�<��;�=���n	��_?�ũ�1X{)<jZ��..PM��Y�WH�S��Ƣݔ27���'��c>4�O�U�g���U�TL�8VV��u-�b�L��u�o�͆+�{&��Wi ��(5�h�拜c�A�ˡ���0FT;!��8����7sr i�O�f	{P6��2z�A�����p��⺎��2h��*�ϜV���:�K���`/zg���`"��A��
���s�����%ȶ@��Բ%�������^ �	�o,-dOd2��%���?�q(|��sݼ�#@�b�=���㳐:+��נC�䋁�(�6&՟Cܐ���R��	�"�< P�fy�5�ࡎ9O���̯��z¾��B�DL��JH��2@I~�k{�.��Fs��4 �g�2��S�|�am�0N�9�d9`���d�	�P�hl^��i���B�e��yS�� �AW���AovT����,��s1(3�%���h7�k���&��n��� ���8�fOC��1O�@֛�>�sg���T�+Bokbh**��E��=���M�O��vR���o�����?>���%�۱�Y���`ڼS�hn�S��˨�3'eލPaZ$V��x�k��\���Ƅ�֍���{}�B�Nl�ٍ���;�ex��*;��7��%��s�[.R�|�A�A��@v�Q���.5��Y>
E4��=�I����V��ʠ��$t������h��A�m� D)u����]�ݜ��o����dn���!�T�!�����,��÷IG,�)�z���6��ho��W���E���=���«��=�+��N@��J[Ѯ?k�B�1�#͍�0v
<���dx�,�h�.rl�)%J����W;�Jz[�H'e+:��8�Cg?��IX�J�T+)1������Y}���"�,P��0�V^ү�rӍ�������k���� z8��$9J�-�ƍ���n�]��: p�1�\5e�w'a�h�
�h�������-y2vgðҖ�FN�	�r9o�ݭ�N�B3��3��?�!T�v��{b�&"9��JP�I�U���VAW1FāI(����Qj���e]r,�Kp���_z�U�Uq2�m943�,u6��81q\���<6Q���ʃдP��x_ؚ*�aQ̺#�����{��`���z����H�{n�~X��I�B���lq���(��0�t��M�_�9TQr��&���(�Se�0�/�f�r�R�d��ІI6RT?S�p�K�������]��^QU!}��w/LK�ma�/cZ�5B��A�G)�0��;��|I�L{�Rԣ�ٷ������^�(���-�%/߹�*�z,/���i�Q�3��w����Sr��Y��z:e�=
ȲZ�65b��T����Q:�>�Ǭ�ۆBI�
XSR�ր{h��~�vC=��'v1��2Ȼ�V�g���1����r/W��a@�F�ݸH�i����[��p	�lOrIj�w��(Tp�zs4�Wo�Y�	b�H2���z�%2��E6�+P�q\��^��g1�彽�$`
�_������S^�!�H�=�g����o#	�jf��U� �\����Al��S� ���+�CӪ�`�ģ^f7�.{Tn�å�j��f�h���O�  ��P����%���N�AK�;��:���mv�����Y<�|:ٴ`�0{��=I���>C�7�rP���b�*6V��q�����kv~����v
�w/R�o�V
����[�\��O� ��1�L�e�?������ a�ѯĔ�$ư9�9��buל�n��@B(�K�����z�J��}5a�b��k^e�5��ϔt�V�Y-�m,M��X_��$��w9�"ѿg��[�h�;��%�^r�pʣ�'��vm{`Ӆ����ӻ��Xt�X����S��u�{H �'�2RO��9�j3��gg	�#����j��	����-��AQ"��z{����;�5�C��6�ʌ1��-9&t�|Ar���C��	v#Qj8�ٕ&R<O��!�{��.X#�!�P=�zK�sjl�d�V�^�u�.�i`�mԑi;��_�H��1�Te�؍��`��`$��;Ἡ푟�����^�XL�"xI[�u&��0���Xv�Z�U��x '������c�{��<�B���HMM�)�k�lN�IG������e�ruYSޙP_��W)��F%�kq��*���}����L��~��V�.�(��`����	�?Ep�]�>�0@�N,!��!�H�zT
%`��~r�1��Y�	k%ߤcwG<k�?J�����PD���nS@Q�;�'Z���N�fᮄ����"-�m�[���V�~�N*׷+��H6#,�0� �C��~����Y�1X�@���:�´P��^�eq'B��Z��D#�K�L
�0�/ay<��E$��=�*�8
�)�<��/��z��L�E��ZS�]l�ı.zR�G#�g����Ҽu���V��	xy��H�E�U̮�nۭ'wG�v� ]���v�Đƃ������\ڴEz �+���'�:�����E�4��B�Y�*S8s��¶�_ԹmmcW�M�&�_�B��)��שl|rϋ%���<�b�1�:+�.oѩ�f:�����Yؤj�nɁ�8��A4!I���m!&r�?�	�z��yV�����u6�-b"�����Ę���8��7����!�.6��7�)H��cl"�͇z#��N��c�9��;n����#�i8��G�	�!�u�	XB�9�5���zi�2X2��x���j����~� ���U�>��;$]�(1~I�YnR{%���q��Nc�x��I<���ص!�88��@
�N�#��J��?E��]� �V�TC�<rm���B���4f8_�$	2�Oi�3,�/�� �7 1��Ap��Ty����*(���m��R%vS��~d�����U���p
W(���!�4 O�)�'�@�0`�5�$>���C��Fb����8r��E���,�O޾�c�����^�o�-��M���3����6��yRB���ӻ����"-��ħ��K���T���O2���j�����QH `1�n�E�����y)����@N�TM�6�p��H=�},G���Ӿ)U6�#O��kzrX�yoh�r�=|C��h��eQ�t�2�}�kl���Y��j<��Vt>9WTʪ��	���.�mT��3�]�����G�P;;�Ϥ}�q�m�*����oo��3l��gw�y,�#�c���c�g��j���
14k�^�g�3sԟ�H���Ť�q����i��s���Ia_���I#�}�ӵ���/�ˢ2ˡJT�>��ۺO�츺
��Z/��-T�^��H��=u���_��* ��$�0����~N@��n���':!��i^�W�b�'	e�q��L���:�2���G��;sG*Q�^i�Po���q|<�k�oAѳ|_� ��@@i ��.���*��iO6L)̔`72�0�����k�S��EDl�N��40����uW�'��i�0ΎnOt�Z�B���Qo��P���d��>��|L�ùGvO��}��Z���U��}�v��j���^|��x�D��L�`ޠ�e������12��3�k<��t߀"�Ob0zo~&m�U!���nI>���K�O�H��̣�
��6W�\�,~6��-�E��?j��>�>7xs��N��D�͡��0�ũ�_�������	,/`jy&v��[�{Ep��5�9_�e�+S膲��o��wl��W��Pۺ��
�N	����с�r�\�\P�����\"��@�������<�'���5��wE��}!3����Z<�X�h̀�)�|y�[>]^��)z )�k�zk���"�]��81��D��%�R��<p��Xd����{�Aں�T�PN�_y]���jr
�=Va4o�{�c�1��lN�Cʣʇz�\F�n�����q~�r�_�W=,��WI���{�2�DFU�9h+d��J6y,�R	R⠈v�ՈAd��mU0*:��ɵ7֓�P��c�D$�p�QN�)�p��E�1��hӧ��r�G��H�yX�W�R�})|9�]�'�S�z�	�"��5�GR4b��Huc|	���u2�v%�P�k�+N�Z+�Ёe�M�7���U�E�it{��$���Y�q:5"H'u���f��t�q��+ޘ���ZK��ZfF#涑EX��I��|ȻX>�k!�*�@*���%*�<�v�6q�1CB�E��r��Yw_%��?��W.Ŋ�b����U9w:����.�FC��	��t�# B[8�m�r�L��U����-��*t}9"���]y�2�'&�>��^)L�x��7�eH���@̉�!H[�0��\R޼=�&'�(1�J"���+�F!��fݫ��<$�������	��5�t"oR'�Cl��(�����R����g��wڸ��K�!]C�������2�%�}�Nf"��O��l�n1|����L��HQ1�x,"�����o�M9��f��	��q���*/z�@��N ��i�3��iFw�I�*`H���I�FX�Z�D2I�����4�����6Cz��Og_�+�ީ^��q:�����?���<�gJK}_4g�xò� yl\���`4��g"hU"Ӳh��_'���1��{S���E�R�K�ErYU`���zK`�Eo;����>��w���ʗ0��ܔ���b���!Qv,5K��`2mJ��m*�k#�B�w�%1/��#|�/w�.��j�Nl���	TN��v��,�.o�_�j���u�C��heM���1�z�D>f�$*k(�Og��FB���5�+ �z/��@��Ҁ��T�F)����._�C��ʈ�c�k�<�JzYkfct�LC���av�ߥ,�X�;���~ �:X�������L�K�$��n��B�Ӱ������[RDtl�8�h��H9�Ӽ��Rh�l��cx����k|�BV����P7B�4�8�d�m��U�Ϯ#�U�e�߀��<�{c�U"�c$���#��h�ɣ*��J�qZ����1�LS�Z�x��8��/�:���#�����C� �CD��s��<�Z�����pr�]����@�W�D���8�qv�г#���b�[Ƕ��Ώ �'&|��\��h�j�w>��ͼ�9U�H*3rDdI��5�O�C�5>[�+���9)���t4�6���%Z�8×����.�h,"8c3�O��ecxK?�&��x��I�����w���7D�����4i5�v���]:�Q����0��v<ꡛ�~�Ap�&jY���uT��3ÔX�i}D�	j�7n���|'�Ԑ��i��G]8�I���}���W�����Agfx�4O�xG#�<��x�2�~g>�u(U:E,j����1�����lġ�[�K�x�v����N�i���EBLBu�,	��(VM��T.*�xw��ųծ�Sǌz�n2����x,���ƦG��)�d�>��������Hs