��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S����%J�b����j`)�u�B2z�l� ���#�p7L�7>J�ו4Ű~;�W�I�]�Ec|f�)s��˓ߑY�u�����|��
)��0fkh˔#�v��b�ɸ�* ���g'�����3�93�w'�%>~07�I�%�E�v�+J���q�[���s"k,B�ɀ(L`C��E��"�*KEBA��y��g���$�~mFy��X���x�,ᾷ71mѡ� �<:% ,I��nu�t`���Om-хb�:ǬۺJ�:��\j8\�(�_�Fq�֫8�+1o��3�p��]��ۄ�Ұ�"e�0����G
lX�y������ͷ�TQ�' z����y��rG�b�Wy����N�
b��W-ro��7yΓ;�e�-Ip����@���Rb4掔2���QH�3�ov��ڑ9[�2�`j��`O^�%�ğ����z���l��.P���m�t�[�J�\�̇��f3�����s�ƛ�@��ѳ��O���E��6*�?��<8�ѹ�r��bk�4��s��M�Сb�`an�&��OL���Q�ť�-9���$�a�[ �R���M(x�MF�5#DdkD����J�A�"Y6�Ȅ����{2�N�d�����Ǒ^5ш�/3����4@�9$1��ֿ�v��e�o��� e�#�$�ߗ��i���0&���!�� vSn�(�w���dC��B�xm�ͬv���Ү֔V�oG�FsT"*I08�aH��r�Y��V	c���������'ȿ�F��+ ��+�=P��e9/"�C��"p����(���&A�DΧ��[���N{o�^��.Z��J�>�v��ݱ���'1�c5ړ�6�G+6T_���oåM�;䕑�ѫk��P���E�+p���2��l�;��SEn�,y�q�i�>:��*0t���̈.�=�>6m�A���툉�n��+ͫ8�q�b1�7���2�kc�;���5����=�k�Sm6S� ���1P��߉3	E�"X]��ib�Y��~�/9�7�J[.�z?��+�/��6!{�~��њ�0�i�[����I޺<a�l�@g�CB�>ݮ$\0�b0ܧ��јG7��b{���|���Ǝ��ܰ�v|Z%xޕ7���ּxШ\��	���i�=�Ф�R�8�Ő�q��x�(iN��=���5hRg�<����]��0)Zj���}�m�&�]�X���=`�r���8�1������z��ʝ3[foe�^��R3O�sǬ��Úd��>���9�a6���,��r�~��c;W�Ap���KZ}s�H�WO>��i�L�>ܶ�ݙ��%���⬅�|85	�A��L-�;~[�>��V�3��7�P]Y�cn$c��%�X��~�/p�x��+���meԬ�I��9�X緲:�hK\�·��Y�W��h6��
J ��v��+8��#zKT|�IU�]�'�TkS�!�C�F�����{� [_&\��>e3��v�8�H��s'P`�͗6�ݻ�L�BOƗ�w29y^�
����<�#�c~ߦ'�����18HA�I��1d(_P����/Gg�8pS6.���g�FY" �Q`	>;ǵ���*�������~���,.x�+�&1�\��ݿ�8	7���h�<�n��H&g}��;��.���F촔A^Wh�7s��X��Cm��a�c��/�r-_�9T��Ru���o����iRF�t����o�#��]O�S=�5d�u @���rH�_W�,y�߇�@� �"h�K�Z��2^P��������	�Hc�q2fe���z�����S�&�U��8�t w�Gz0�b��
��o���\�ɚ��!�WN���Lt�U���$P8�[��\�S��35��F���X�1��)�X�>�����^M�����+Ȱcx��z�����?:D�I)�6�m?��O�2�����0��bν�_�17�b�M�̄�����MP��\oQ�0z�������Euv(�P�����dKoHr��{& �Mv��� (�p�"��=槏�~N��$��_e�^�,,�
u:���O1.��w������L�T�����X��t�/���]3c�)��qNv���>��mW!�.1�r ޅ�7rV�4�3�X���&���S�v1��h�rMO���)�"#�m��k�(�/l��@կ�l�c��ܲ c�1�=-��&$�]!�ms����~ �Zb	��Y�ݕn�-�
EĔ}�U4�áɵ_�Wz)��I���A�g.B=�݁����0y�O�І��'?͖6��U����>�jX4.�͜��E{��[FK�Q���@X��y�L�gqY��PԻ�����?cI�u�nh�a�@-K+�1I�ˢP:.�bV`o�5kQ����ej���e�R��O�4�U�H�9��m ��L�00<��JAS�����Y��΀BG��K�ڃN.��Y)�3�4#�q*�-��$dT!�L]��%]�{τqQ*D��OZtO"��:V%���� (iK=6�]��r��*Kl���Q�i_�=���t�2�]>�Exp(W��pt���;�n���!���YS&䉟�����Ｃ�P����NR:v�z�-���8)�F�=��+�y/B�������0�rX2����E1%Y�l4F����� '�l8F�j;뵻8�9	��|<s}&����h8���ߋg��d�aE<t~���2_�*c�:0�>��4s��pOs�|����]��}Z�Y�U���wZ��r�"ʪ&��qc]�-N�/t�0�F|&�L=g���?Bv�;Q�L��?0������*/��z��YX���! s��m���l����I��T_�M�����O���[�	��[�N�-�|�En����P����#��XKN �'̚y6F�ݧ'�:3�[�u
�J���"�]�[0�80}�þ;�
Ix���gA~c��ޟ��yo0���fi՞s���l���h�?���Ɍ�Q
9��� o`?ZQGi����HhT�z2|�	UP(VzRc4��߃ߔ���]\��N��y]E��U��i��%���QNZD�����o1'}�_����}ɤh����38�e;�R���y~	���XL3u]C	<�W����a:��o�~[�#+��NB&��-6Ι���e�Q	����,"��P>��� �a\�;X��Yw㻀v;%+���Z��J�?L��� w�<��&��Ύ���s��{�s��BT3<��h�Q��"SJ��"��g[�hS��_��ݺ���a��{Qi����XГC�ra����Nr-K;�do�|���ˏx�F�/�
�=Q0+F�3Ґo� ��E��}ޥ9(܎���JIAb�3��Q4gݲ�G[�R�Y2/�V�'H� YZw>y)o;���|�M|Z�d�g��fU�|3��4��ｇ?��G%��m���j4uj� к��x6�����@��ܹ˹U���,�g�����I��n_i�tl�@��x�� w|:�y��[\����� �62t�����^+#��d��[8 �I�����r�V;�ƭ!�-gQ�;k�F��ލ��HY�A�q�[���,y0K��-C4�g�-^eQ:�^z��b���֖{� �e���Ґ5��_�s�6���m �=��c�ĸPb�'�Ǻi�{��>L.X@�0�8E��
}f��b�-�������_y�|k]�ڵp���3��J�ψv�`�R�!v�f���T�;YJܡu���������'�=��.��N���{=L��I��R���Wl)�[���Z���DLd@)�G'I*��2�	y�c���1��)k�_L]�ч5P#J�EkޠB|�+�(ů�%<)v�Y���3~LǨ*�0�g��%2�m�"�`R�M
��\�5j��]��X�Q����U���9Ǘ�.s38+M6�F����5��'H_ q����D�S�X�����k�	�+�j��٪?���Rs��wg�������A�L>P�wvOuY�~ht�U"���n�x���D�mz��I���byZ��X�T Moh�!2��v]�|�SN�5���pR��Ο�|�Tk�R(�?O�o�[+$y)2-��AGǿE}7�̦�s��y�a5�j\Q��
����\o6U���J)���2{��7%G�V��@��~�zν��]��s\��Ǘ���������������ZJ5���7[y����,��ouA��b,ZTHV����E��sқ�x�D�����k����?�S��|#��E�@�&AL�T�F[������|��""��y�D"K@Am���H]ڢ�ٮĥX�F|�\�ȴ��É廵��ZY��UJ:���~�i�p��I�G�Lx�|ϯ$]�2�Z��*�pn{#�cg��"��w?��s�=�x_�3؉y����}R��U�8%�3�Z[�N��hn���j�E݀���������K��8h�2,T��e��<<��܋�Ĭ�5����4��Kٌ9S��~���OX���UZ���׽:`e��E��qv�[�FG�n:����4�u���n�ig������S5���n'���P�Y��ms�-��!�D�e���.	xNZ�kĕ�k �'�xAVђ�J,�ϫA^��� ���$�1�MS��A�PKL�%�ߜ�0X�v/���9��	�B6�dR��g �8ᚺ�'>�^"�B�=��v쯞 G/T�ݢpt���8������ϧ%�M��\l a����g�_ac��]`����������>	�X�N3��ev|��=2BT>(K�[|5|5Z]��G;��-F��I�����@fEV�h'45!i��񇑛��q���J#��<��nTЪ;��`��a��,��g���h����,LQ�ڛ�{<�bL�'R�cp�I�����oZP�q�$۵�k]T���z�����dl������H�"�*k�n�E��G�F�a�9�NZ|yvFT�R"
D�UD�~G��({N�S��,�f�4��L�l���}�UQl�V\&f��ku�W�H.��_�e�]g�ԻY������9�ڎ3�`EoR�#$���?�e�d�
�L�"Y�r��O7m� ��D��"{�i'e���n2���W?���P�#*#z&F�!�,�[@��;N>���ͧ��Y$�I�c�������̠ٳ����t�ޯѮ��_f�̜S'�/7� �|ޅ]Q�ӈ�HD�')F[nµ�� ���2�Xʥ1f]�	M[48Ҕ�J9=LH�~�x�d�S������V}����D�ZfS�V&pk��e�{�R0��?��Q�̦�P(<N ����r�����[v� �h����ƀ�:KR���:���ޡd��b�Z�'o��7���DZw�\8�C��L>���C��� Ľ���[��j�������&��P�a��j\S��?��&;�>X�H�-A�LW���u��}��"�Vɰ!��ݿt
w�n#���C����?�3�)j�I(<T�n��ڇ1��n�.	t 	�f_����D���.�Vr1�e�yf��=��{BP-�������h����l�EO'�aB�Ќw�ڭ-�]#��'�������WV��)vj�V&�h��t�	VQ�"n1��yS�4��<���a�wkԮ9�)��S)�	�hX�E��)1��PFD�yg����T��9��Gi5��ߌ\��Tk�2��ϑ:�w  ��}�^�C��&2v��R.�i�6� ����a�U1��Vx �f�9��P�BM+�ɓe��zJ�ؕ� 9�08�;��'��
��X�J��@R�j�u�.G�2����@�c��O�h�����Cǎi)n	-`��ńx�������Vn�L��Z\���(�hEUW6���B3�)�����`�/E�g�=�����f�rG��I�M��hm�7#!$"e!Tf���Z��B�`X]q�bw����15l$�wy]I�^K�Ԁ�U=�(���D[�����'\��(�� �)�����u��>���n�Hxo����Sލ�����h�ׄ������B���Z6ߞ�c+P�2��q�GҘ%Yt��>5����Fwh[d<+��-���C|���'��x�=��e.�ͱ���%/�����E�~�(h
�Ml
i�;�"��X�σn�+�o�f3�ud��ˏ���eA!悔�,¨9a��*�L�W�Hhf�l�=^���j�a���l�h=)�}��BC6	'������[�=O���`K��VW�!5��Jg ��`�CE

��U!��B�~�W	�|�l��g7p��.y_/��e*	.�͏�
x��q]��Z>���2��T��b{����9:o����XW���o`��Dܿ�cJ/l�a��{[
�O�F�b�W�0Hl��X4`�!���c3�|fZDPr��m��x��7��@^�(��[���Sy�M~�'���W��Bu^����v�y
�:�r;蒩��ߡ�L��,ZPƔ�6�C��,,q�y���]9�w��\R$�U�a�jŖ�!���2���Y7hoGog�{O�^*�Ow5ī�.˷J)^�� ��\�m|�"ıC�C!=���r��ŀ�L�����6�\��Rso�xg`����D�<�
\�I���fD���
p�{����h����8|P�UY���:�
��A#i�d\x��]m|cb5)�k���#u���z�+M�cG���y�C�G���n�v����!\�w���S��\|f�8�%�e��W9ë	�L����k�^���c,~���Cƪ��cD�&=jG.i[L)ׄ���<^b� �Y�D��>U}��c,�Z���D��L��f+���pO�i���KE�{H���4�.�M�ke6��c�LC���|?�k�V�D���k���4p�P���w��*��c��CV���ϑ^NT��6)����+G-sw�(��̺��ïb�i	��6"�(c���5�J<��_I=ې�2!�&��>HEK����k�()
lc��ؽ��>��%
���/�=$�%!J}_R-�߶�e�m��G�ہ��/�nɲ�J��t�ۡ��������؂�6�,T�`L�n�ʴ��L?�p2ް���j��U��y�1�5EU��V�¼��=�q	D�JJe�� �����F�V��~bX6�!���R�h���} �!��:���N�&|./��ռy=��"~��yp��4��I��jsW�����BuiF͖~#�ZBJ��c5�|���C-Y�R���8 �����#���x��׺�l5J �ɖ����_-!�o&<7�&��%;��\��<Ōxa�� ���:-<�57g�Wī7t��N���������W2R�����;��e��-��0ZN&&d��0�^H?�A�x�|+��!8�	`�,�k����Vܣn[^�U���U�lѱ��q���c8��Z��=�J�+z�a��]�y>)7���<��цʻm!`�n�^+>>jL�%vE�lyƉ]y���>�s1�R�x���p���v��u,�l�:��!��� A3G�l�:�w܇;5ʺ�)�V��ŻZb�j���_���a6����aQs�����(0r6��X�B�4ŗ�ڈ�=�[L4P��`:==�<d4�H��hS������~�Y�,�ƗXn���^��Q�$�=Th��E #��˼�I���g�A;�c���>� ��CEW)pBw�x��O/����ޚ��p��o��m�|���A,׽� �w���Osϗ3]9�d�\`Q�~>��|3��5��z/�ʱ���Ɨz/�m#��BN�5ӢcZ���6�1�G`m1H���"Za\ʩ \.����=�\����"���Y��h錠Y;ݴ�/W�}�-��+?�!,�'8�AGP���'KQk�p�S�8sTo|�
�2�o6ӦU>���@����	�	ò��;�E 
E��zш�|�=YT���n�]d[X��iR(|g���p	}/���S�ܼۃn ?�0Z���|.���Ǟ�s���U�G��T4~n`T����ׂ0�|>��@�J��c�}��OBn������5�_�e[�H��ђ�Yx�dX��ty��z.`��i�"�<��^q�!�`&��{�=ճ&,<��F�3VR���}�6�1�2�>��ٯ�����7��Z�6�kn��rY��ڍ�ځ͟C������T�a�b0K���$q���E�8�3��{m�#^^�� �T��d���ğ�f�k���(ܵp\�n�P@���,�XU�؂�+����26 �Z�ނ{-81�p�"�H�Y���6N��I�r�-����a�w �PhmG �C,���d+]���0���=jM�#����$����@"��NΔ��
f.P|,�f�t�g��K�����o��� m�LC^�]�}�E#�#wb�mk�"֎s��N�U�|+����Ճ\A�pͥO�k�ASJ���T�j��/���;Zx�[ߋ�.�Ԓe�v����w�.���� ��0�挓�Y�&HߘCa����� x�r��cP���`���������"vt�v�w�J:Z+|?�Wc�1�QQǽ��v�L��)�!V���&{�#f"1V�M�ܡv�fQ
�/�{�Φ����U�����s-�c'�.�X�.Q�K"Jz7r��+-�+ll���c��wRA���j<�s�}{�_S�t\i����/�<|k/�ۦ�o�EW�6�d������&cxBn������ｊ��!�|r�E��ZQ͵$끩�EV���� �"���;������2���=�p�φ�*i�؛g����;-��0�����97k9�uQ�g)3�d���Lѻ��,�A� "�21��|t�K=D�q��A�ࢨNo͟�0HN�����g���B��F��F~kU�ؠj�ڌ���3����^���Yu��]4^7ay�3�o�,=���#��$Rɷ��Y��� ���{�ZH?M�(BpP��!��7t��$��_����2>'AҬF3�f>&T�Y���fq��U�����A��3�Is���gݘ�Nv�ncYJ����ۈ���G���Ƌ���LO0ی^�����f�j���*�'�B���Y��f��3I7>#2Αא���^�Ĩ@�L$�ה�x����z�O�i-�S�Ü�Ij˱!����Q
�'�;⒂�A�iL���+�~�v�$d��̅�)h$���B�Fл֌4;�e ;���"=�����o�'��K��Sݻ`�!ޠ�����3Z�J�0��f7�x9u�
������*���>_G�ўA:��
[!�-L�ܳ�喻b�yB���j�Sk�G	��K�&�(V��4kK�ߊ�/��_�s�C[����GEo[�^vS'W!fV�>�d��-��WqЎ�q.���� P
����|`Ϲ�Cɣ�L�Pc��~�Q�'��b���W;_զ��K�K��D�L��`�PZy� zZc�*bxSy���:R_��k��=�����t[��fz�Hi��JV��ľ��K+os��Z���6�����nqj����7/�ˌ+b�8*�0�ivo�+�d�.&�����?�XFR�<>�N oC��\|]�@��]yu$��;��xYð��Q�� � �.� �^�6�5r��Q�@���3��co[	Wg��|-�@	X��_�5:��ce]�w��F�R<�k��d�	]"DgQ=���a�~0���7��_�

�����2�i�NB-��v2榣�q�� �vw
�9�[����Q|���_�O�b4o��2aR}��K:B�!$2��?(ʻD�A"�*�?�,t>�8%��]��b��30�d�}�и��s�TC�ڷ�Z�G	;\:��6$��'eh;�W_��:��$��?���*h��t���M�	W���<�3 �Vj��)}��&��=���,
)oS�}���`G�;��0^#�����:��7��CB�n��=�UI��?��UǢ�F��:L9�?�#ͣ��%�``L��v�,s.Q�2��lj�Ss�l'	��-��z8��ۖ�u���P�E��X�� ���=^�i�)��e�X�@��?�bcxG���c�T��.M;�|s��{�[%ŝ^dtZ�cn���L{��21p2�y~��|l�
���!��e��	���6f_��6�K8��1�	q���� 7*��$'Q%C�)6@q�g����M����2���5I�D�����&�ZyX}(/T9'^qp�I�X�j๵�rS�L�����y
��u�Ig!(Aq�#�'"��`�#_���o2�@�'ͬ<�&��D�w��ʜ�X&�'x�� r[�f}��<��RQ�L'	J)q�V/��3� GY�ά�ߥ�(b���R���y�t�V��5��ĳY��[��@;)]��(��g�7m�q]p���5v�XBuʞ�g����d�9���~�̛����i!��='1Uy�_�Ob|��Ŷ%N�qs��: *��6%p��	�5��4D�S���%��@��Bma(R����nzگa��=ϴ��X�(����
�㽆���2��ɋSm4�+4�i�q�sn��h�c*�b��Ԓk�����Xo�o��n��4��D�"t�6"۽y��zV���Ξ��<WɯX�g���_��������7����$uݣ��H�_�՜��	0>ȧdUg#��N�sb�M����)n'� �)��u��{�t�JYuH/�Ix��6	:0O�8���h�4�[��O�J�o�Y�:Omҏ_���w �^���n���=ȧ�!����2������*grxG�/��F���N����}5�F|����u���ΩK�E��ϲj��B\0�!��@kb���zeC�t��f� �4�(��w��/��;��ݥ�R�~$h�X/������y��IW4H�7�l�s�}�^�J����#�s�қ��tjH��d*Q���e4�+/�������܍_n��p���W��=��t#�98M���mԱE�x��������&�g�d�𹻲�ޫ�T�w�.�	Ӂ�S���G8x��ֱd�%~�=�� ec�t��Ճ)cښ{�݆k��,� �B�dO����+��(��D�
��h	m�#v~�H��T���[�}�K��Ȕ��S����F�[�3}�Nr�r����5�9��ow����oР���q�=�<p4�NV�����=��O�����4���6i���2{HE�Z���@w`clM�̵���f7q�� -�8����ُ���ԋ�����2��!o>��m.����!�:]�p�]���������l�9���*�;�+(�0�Ǵ�g��%�;��q� �w��m\��/m��A��'_�3����H4�'���FU&�ͱ�sR�eY۬���m�l�����K~�W*g�$��j�N6������₇��A��n����<���H�op`-�7�1��\���SM@+�ˉKŶ>�:b��["�̐VZn�|z�%/o�z�-|$��h`�]�R��0��|^���=sl:9QXpͅ"�F6Ē��>�����/.���(9A�X�ɚ��Ś�E���)�a�Ώ,a
�N�*<�uN��?�`�"�
�4�7�`�V>�oh��l��tb`����A:�s&�Y������ۇ��3��/�5rx��`>B�?��0��^�CC{�~����3)��ӌ��M�����m�|X}�$M�@��a��L�Gy>�H@�w�;�-W�N=E%�Grp>Oq�n����(F���uB�m8
���y�J#ߔ1S|H�}JBL�hE,�Dd�)~(y�"�%���O��Zs*GlÀ�#ݴR7�ƨV�U����¿���DE�J�-�t��lw��T�]��Z��3��@�шOȱ�[+��KKVR�p�r��_�>�>�9��c[�c��(��X=�\;�,�a�.��e=�g�G\J1��M� ` 9Ʉ�
�HiҲؑ��V�-(�n.Dl�8��g�1m�T%,9k��o��.����8��0��y� nQ9P5��+Y�����F��-rL�A��KR!�Evn����lp9�F��`�"Ou���'x[c��:S?SFp
Zn��-��G��0�nm�D�EG��:���6���d��)'�.�.BZ �&��]��skYx
t�����xG��v�]؃~�*��F��\z
t{�37�_�p�I�|�G�+;�1�)�Q�;�P`��l�W*mm����A[��]i���X����?"i������� W�9 槃�?��냚�ջ��6:9%s���!���.�a�\v�`��:~6>_�G�B�>A�<��M<������^	"�Hev �X���M���`�3�WoK?� �w+񵅇�7,�r��JĤ��NEl߆D��.����W����|�P�GX
�Jg8�N[�8�D{��������zB�?$�٤
�g�}[3��U`��?�o�Y�.��Q����&�66� ���g��N��ˁ-�¸�5��w�1�X�Ի�Z�04���Y�3�;ҷ�h�9�g�c��5zϿH2�zvp9����΍8���7��̵1Z?��ck��7���b���`�9�3?��P���΅1��I�åd��蕃��
����O� ������6&�	K;�iB����5w9�"�{s4�"#��%���^6c��nx�������9���t��8
�����B9y��V2�M���R*�YFپ�\��ӻ
u[�/��h&*n$�a������ɾ�������sM ��|=�_�V