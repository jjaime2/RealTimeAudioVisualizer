-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mnqsFGirhrESPwxoPybzc/hD/fNBu90WMoDvXqfirlc1AKO8qAxcwyVJ99tqd26hJxRNnQ4c/icw
Sfjdt1jtU+tStE4gtUKARrUEy+F9GWU9NNgC6S2HN8J/TlNzbdNtcVTKpYv9hLF1Wts5RYKSJnx2
Wxod9enjSu/purYu+Vn3yuFD9KKNHzacscv1IKOJbZjUqjS/+JgQNsIrxW/YO2wQBYNGa/nXU08E
UZpmZp20Ro/k7aPcwUJRsd4wZOnzK8zDe94LEtsZa2zTZQyapoqaY2wswQScSKaWgORrN4s8/qQM
scGYwUIINV0b8QTuZxxQmEZo8Il2mp78Ru422A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4976)
`protect data_block
ScY+rnkRM/ERqIrut/XfjYF0oVmL3bjCUoW/OqNIi9RsR9tFDgbdgjIvI/99ldxqjMPvldtAZYYK
fM3ltQ80P42/ZusUN2jADGxb2WjH1TI253GxaPfEq99/cSWqFoBZspUa/5I71btLYAkCnZMpUezR
qpYl7pYlToVnw+1FSX5ZxyCEHdEv6sZ7PFfmocqfJGIQjKLik5xrHo7+DlZKXdJXWVo0GdRflQOF
YGnorjrvaibkT+X2TbLx6weJImDwnzLAxtHEDNyc+gf6CAXA3s+HH5JUTlhGR26Ew2DsWtkhksCR
G1D6eKO1Pdw1ljtGKlmsYsXNo1l5Jj2uNx6BXKxob4l1zOdYZsSsefjF+MxljlLm9Pcnhyl0EJ9Z
Y+gg7b0/9HGrNfMGZxKFW3BBWipVNE0Z9bnnuBebdJhkfXXTIv/3lo0z9TQbK9wy5r7CTrxVJMOX
BGRDE+wzLkZGk+xAfDjJuTP9HAEXWVJJUt1a01QqROn7u+5K6B7/iKHRhilgKQKsiH2Cs1V3Y0Q+
O7BNPsh16PAjkWn1Drq6kXfaW7HuM1biVt2IaEbiYAdWeNQ6KiVzsbi9JknRLZb/c5o7xal+lNj9
q8bWJPZm7Rnp3ME1yqbvngDKPHIrQCTAoulFI/sPMFHv5QLpPXceeYbgo/bgSnR+k/Fo7JIRMmeH
e4TqSUoPZG0Wx7UUrN7dR208aj26hTc6Lkyw1fuEfbpTYYqGO1H1Eny2cHcZEeHzcPpClRYYVn8f
tA1jypFnFjW9L6rMAUTNj2yU3VZXtBKKoAJqZGNtgS2su1c8i1NAD3qW/a+kl1duTbse4HxYcWRM
uPmxR6x11PZn9sXinkt4aGi9F4Artu/hBcWHM+I6kxVrJ6F+OiFgvs/1Us3E3VYHJPNJq6t6dDsN
UkfQ/1X9AQsEOfp0WfeBa1cci94Mr0StIXVsiQ696RC7cpSHenzHveM+hZswpZDo27auzBE2d5Xf
ufBojrA6dPJx6SKFnh3Bw3NlPv6FSFJmZwnZT9RhGhhE3EqEs/HbVRrUxWlL0zZ++HmjuRND/6LA
3C3o8UU3clwE8UMofz0ct0wuX9HzdVUga4MF7KoeccdN5cj/v6bAeZiuTYA1DjgtrBkoT0bHgwr+
aDOV5vPeqExb+psU6KbfovaHK+ZdS8glKtF1SnqvUUeURGmsg8UzdFXYU4JsND7Nw1Up9+vHsOhb
2cgQ/Uvhy0/d4Ja2/KA/2uwU0mIEw/SBBp0yLEei/1tDt4SHRKCN3RPZW85DIaySvsgpnNvqSzb3
yXOFcfGVRJDH4rR6y+nxbFXYff4Ne0pb08t3iRnBghZ4ixMeS25EEgxNWCfR3ReRdGrjkBTfsghv
wLevpQFF/ZyUAJbNrlv7AL2wybOr1jW7z9oo3jFs3MeiUrzMVxSORoWXeB6U/5lC2bs30e6GXkEE
rFC8ypOaOnU735CCtXv2k9VgBeOSdTRnTODzK0WjDoOLKzunCDjdfoQY2+fgAm7bkmcXBHhhdYuZ
Nr8aaFb4NI48KtJ1RwPXCXJjyr0e4169vN+mtSuOuDU/3IyTC8aN1FCscGqEVsZpPn5V/r0Ga6CD
pBKSaxwQ2jaG0fCO2DiyrcJLM3EvTIhv7CYyGPxz+Ml6v1ZkzjXrCroZ9CTJzaDr2u38EEhJPMvU
fJGt7vIv/FQldamNAKA5OsHllXdRpDvekOQZDPBfTx3mVTJ68dFvUTcpG1aakxV3e2qSIK3Pwf0q
/xLkbIUwjKZyjqSMtl3jCDoLzgoH/oCH2I2OohJ23KCRaue9dZYA8gZTo4D0/dWUYWKwgNHDNfqf
P6pW+Gck4iHwJCzVC7aHDH6umnnt/8ZiGO+5Z6USyOCdDpY902LisgTlu3T5sZ4DZhGFfLtoY5Dt
Mfx2bj6kcOx7abJOwybK6l0DhrzdLg4weRTQSTSatjv4EI7qqiqk7DJTJfvFAntcZQ40YnY7fDAr
q+bmKf0CcpVYaElmO5Zpsn3Gste7toOOqoJav0++Jhi58k14DfMUeQpT7XPJqGuTEyjWs39+ltpE
MKYhFTflQzQjykQQlor8SJFlRt2TkRto8zxJQI2xgN1BT5OQeD39QjeOaRZTPDCo+35fYwbF4pKF
h4H9oCPIy3sppYdez8jpJcKyrI8IesLHhUY9bCfgZQV4c5um1bnSYdiudpX/Mz25bgHemczf9AGc
HJ50yyXVYTLjaNQg3eMbrZItwZAeC/HSiRlzNMsQWq5I7bixZrcW1NooVWilvocryZ5CrExfozoP
fgY228Bb7Rn8D7ilBUYa3EKjwF+QSVYpWWc8SuII3SMdQvtRD0KqAcHjPFkQcgUnwZNmwqeYqjnP
q+5pDDjTI1/OsBFPD25eVJnsKMt4r84VWEYnPnvv4FV1j3+YWLED/HwqLVNfqwROUVMaubf7Fe5q
KiyMtURV9h+iUXVGr5pJvUrNpgsxN53u9TU4I+4nDoQRN8ptAEaLS0U1hAPbWbdPgnDEbJq/Iyz6
ZmewVl0IQup9Mosj7I8VyD+t0Ix3GCQYmU7zaw4NJW3dB2Vmk2dO8WetxiAnaHE3AXDPSYxpVvDZ
hLWqs3Ut03JfLCelv7oSMlbTqG+9Tx3UzT/l4rm1ziwRzqSwEGjKaMf3sUTlR572TJkY4/Zx97h9
OPS/S0IgHSGjHUqullBc3HqpDoHCJ3cC6+xzO+aXZWISnT/A8VFc0wDQIPwvJYf3Bb9/oMoJnMPs
B9QsLX13aBYJCQBRxQHQSPTOcyxxOXZo210TZ3hn0G08JoYD2cXRJbsr/Xg1uN9lsVamDHVMFZDp
BS7BSCkJ+4d6a+2iAInWLg2bLze+BT5ESC5ktp8YHG5Mo+m2V7QqEqa+nQ1YLiuUsGttQLBOD7ox
Rf5y0Tz5Kga60Lq4YthvtxJD37dclOro4a1cjABcDvzNpIH1edvORnxUm1Wlvf3BR9baohFTOhIn
MNCKDuhPgp7DY2PXOSc1pR9BxdT+Neg1UapVjo1sH1aBWzluo7McLlk7gWI85x9sNE2sml1a8hxD
HmaIDY/2SSpxiOpx7kzPXsTdhoAHOlCOyvNcfQO85zpw0jHXgMtR/vEw78xZaWoOItOrc77xiGer
SZA1fk64oFpxDERuTXiWoQfdXf2aYntfoWeXomKljXyh/c/Dv71ZEvcTsonhcLMjBQaz8lIGeMVN
wmoXZgTrVahf3scVIFJl6Q5BrhUMhJZgMuyUN+7k/CpTqJo8P1SEXXa9wr5kwMnRwri0umv+skTk
JOtV3UmRSVcF0s9+HA1HSP4O5i/zifw9hlW+jgK9eWB72wAHqvLvTgfo7CoCjC72ddvhvcgC9RSY
QxTqpB14AE6yrR6prAWzlYYgxdjCgGHpXDFopxrFEBWT15/yRTw14CwO5QDDdIE/WuM+0bSG8K5s
U0P74PjFHZMuq43Wc5SYa2zhDue5yMfF+DPfKXyWTkSojw7gEyUeklDBfi62RHQwfbQtOrwIVz42
cXVCf2MP4dAcgLZ4wXSAMFhkOoNavGrLo7lYIReq66k02nVte+ApzNarNOxbY7deCcWzCDeqVO98
b2jfWQP3ZUz8cpFRXkKoQLWq5E/dk5vyK331ct4G5PnX+tbnDIGsbAq+f96sb2g72ym3HkkvHDPs
Zg4CJNFWCc6GJrG/WOxOKqZAvTwSfTHp1Rhr8eEdpGC4KmThZtBzI9OdqBP+WZUcSBITeZPglKY1
pknlQRgV5eN5rtGqVQ9lreUIXLYtKCqdnhGz3s7AbUPSDFB2UrCbb5QDtDU29BFD/u1lsKR9z62r
pEpD4lyJWlG1fQxicOAWGYQI9hVWCUJyEnGd+WNp2EmA8fbG4d+mt4fAVBVXco78BURx+aJBExoT
ullM7BA4C9gUcxAayrEXJyrVSA5aZ/vdYZStNcdWavdW1D4d4wQmgHX5pTOltIEzolX12EfUcrjx
7QCCFH4s8crco0btrOZ4YNvFeouKezAlIJfqe+jmf3JPbk0bLq+bjGyu5J3yfMUwVJ7BQxKsSWyE
D7NZUInQKU5K2xUyDxk4A55xBmJEX0Q/91GFF1MB11JdxoO8tsXQfqbZHZkAReiZMWGoOPEqLjH1
01uFZrYoo6B9V8ngLEeDhJw8T6/MPszYGa7YDnDKf9fDPNFYt6139EC5zuV0nEbLRSEWaIx0QKKY
uFnQq4ujqPwBEKoTCUMmCM2I9uzxizdVTFXnpkmrVriZ3L7iOp8as9RpqIasONbkFRnzp/2pnw+m
PSZZ0hxutzDnqk24RnpDk6PNgk2x4dkdPDoBPprLIdBpYIYuanAqahp2kHHMZxeo5rbVKL3TPLl0
p9NoedfmKvEGdDLyPj50GUkbeLnXf7YFpcjK3lsWIZ9hWFwFq5zSc3Vg++KCoht+cYOVJv5fKm65
/YGTxw3vRuSIbgjOSKM+TLP5mRlNLW62EL3qG5QQFaFYIbpU8cZ7AFGTXns9fY2xcMySU5nMc6C6
wMbZUEJrvBVzbdl9koZjHeHbsL0XXeuabiAMtTgT/MDw9XLxi49hYCVAPy5qfUeTnMt9DXOyW3ej
hqLFnBT/G9O1Y2H/ZtxuutJr1+T5lN0HKr8pMko4CE34+l0Ke3E5YyhHU9sIgAheBYn4k400aAq9
TZCTr/Ruy7rLMZp0j2ab1+PY5z8jyX7w1BwAOUA5bk5Ky9fYzJp1Eg4Km1NvA9XhYxgjYD5O0qL9
s9O3AvHVu5GhFskYM7TcL3qMg3YUdUDAxtnrstBiXPNPtFW5UZyeBXfjJVJ7jAlkLqTHokP4G1Z7
aTNjo2meNlmwVQswde/yBea/X6E6Nq6tNwr6zjNedxVPkKrtGYtf4223rDg0zxgW/HCCvXQZdQvX
qrt8VB02viVZdfsVPVtsp0Ttet4g4SlUFgVJ4F0Gq3vlEaEm98qPMCsQCsgLNGKFFrMxlGE7SBA5
knJ+VyXjgCd6CJT5Ob/ANdojaQo08s2RGfhrokGU4eSCkNXDTz8ZWdz1Iu2nEGiltAoUOprW9Nff
rqOiz3+/uSwJAN0r2kT+09G8k68NkoQ6yUi6PQ3QtT3h9kDBPJeSbMFXrLFgrqUYeqOMw5GIQtio
DiBleP8NKfBLVPfLFIECpmdxKnwuyPN00cdmDNUJc7n499Cwgx3HjMn2AexrQhqjkkR4nw0aIc9f
LkA4gpFQsC+RPmgUOD0AVTVvvCP2egJqwdqRNnIcOTw+1ljZjaKBq+BSfoCULOiCGIkmA7wu70aE
ILKpQ5iDT9CSEGFFrEI7SzvhivGyAjIGd7Knp/9l+n52JOn3CEcNNtERsZLox0Mt4JCUGX3bM5QD
wJMHz5dIqx0FbO7vLsFA43Uh9/i9h7TrQ+aSfRNPJCKDclfG1H4nQK0luse1q4+6lI0LNs2cbg63
u+OaUXAT9V0wTBc0OjVCmnJ/bwy9xWi7ncITfRkJupgISNPwpC6uuMK+cdIyq/BnUEZ+HBWJvLit
HYNbCPMpXKCd2YGDryg9F2l+bqcQ/W1Po20hnlcyQCwcbu3tQz2EMc9RrOLJoNEUOsl9GM3O6rnU
WeUnxUk4jGqOQ0FZeyCi8wlLMQnkByL60OMEooHISXaagnJVEOlBV1es1+o1IWJfg9V8DTQ2Qjb/
xhEc4Vz44OYY1jjZ8sMrvQbpn4MIFxqFRnzs7e59FqbvwUm4CATPiWKCLfhnpAGsHQERKAuL0n16
QQ9br18WTTC2lKNnXbfYiFzC6oCkBlrm9bESi9ZQGF7mFltjCA+erbn6rTX9SU3WooA8OuVU6bQb
O/hsMu6FHbEx795LV025B2iyxFlA4hwJshgD2A0qgEN9kntxY9sahKlRdMMBAzQIVyGra/FkyC3i
0HmWFX0ZeVLsjuL2Fn5qoVWhnogcb1sUDQfc7+mBYrsstNks+FixbK3fE7yjdM0tcAUBF/xdpRR7
DbiU1V/Qjurm+Tmx1rRXdhf2BKcvvDS+kcyJ2zdZredQrW0K/DD7i/Kkzt0VX/bfe0EeosCwAMUr
FTfUknYIZTWmzis0YCtcs7zM2QUcQEVIWKsDIBzAaMDmyj4bS+lYz4tS9cPjD8oGGYGlPZZhu18G
8BZYk975njS7mJey3SZShrKPZ7GNB5nPfzeGiyzoxjzMCSqLOhg3PzdjFovCV9uplUtI657FhPwB
tcv4KqeQhIgO2ATZQVYMwaoQcNNh/l4l2PeUc5wA8dkis8KZSnmhi+jQTqJ7ukMkCwblGFAu/nHm
pAjkDXGa2uOkINiLQBROfOjPF7QxJtRH8QaVK7pToH+f2LlMBGzm/LBP2CxMQUORs8RSny9IAyko
OTw+I4+gmCRh8o3gjbJuWoT6H4FxyKrMdei6SN90ho3FkSa91J3yxCs8lC9GjN6tpfLcUvh6fwqg
lwmpdRCEcV2Ivhytu5FuFL3P9BKGfoE/2xlEnabPYiyAs8RWLCgeLi//NMs9mA/tY7EVgwRbcRgi
ovpIVNjP17vjUWem+SxjByuRacBShjQHIq2FCQ4J7wBh/5CUmy/N84kqjTfdcT+pIEVDRy/kdeqH
kjr8xGOaEz8Kgfw/qi4UekvnNrx3/b7qLsCq+cYNelKt/4Js+cx3iUbZNyKrqgPABhXvUkAqsYUz
7Su6I071O3PfiO2wHp705dA=
`protect end_protected
