��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E�ﻏ��Aގ�~ބq\�l�1�4QQB��t�
�_�㬃1Iw�$�=�\�:�}Օqգ�$�ZB�h��NS%`2#r�e��c��B��FJ�CH"!��G�D�}��za�����<vri���Q-	�d�!�s��'�*�bOL qls	��{UŚ<R1l̬9��)��P)ۇR�	��� ���n�5p;D"���mZI�6gT��z�6�WLg45��sͼ׬��*�u���S�!kj/��v�!h̓v�ӣ���?W2w�1��i��B�ћ�����fñ�uCnԯ��&�z���)�?p�e�9F�����x���K�>����g��?�L����&�"���z]�%�;�9w�;\��|.E���z;�E�ɸ���1���Ǟ����965u'��<2��o9P�åg�Q�&���:�~��o|�ٺyJ'qF��W����\Gq��D��S�E�]]Cn�K�2��$M��f��5<�Z����)����Q�����+d�����5�/O7��{3*B�|��C��X�m�.lR���9�S@�Hk�`��)�n)[�X]_r����´bx�!�
���k�g�$I\s \��3�hĒu��͉lr��W!1dS���D�!I��4����5*ސ��#��NRۊ`���s��/3)��Q�W	h2��yI{�+tJ�Z�p?�� �)��BY%1�{(aC-��8QTI�˜4���j���ϡ�%U`�G��3��,����*�5S 齏��@�#�h�NJ|:j�y�i8��k֌c�A�e�l��}̄I�$���Q��!��E�"�WW�s��u��|œ�?X����U����N�oL=bBC�_.x��������5	��VE�Z��$~P� �i�^g~�e��~O�K�#���<��R�j|�ւ���v����y�o��G��;�o�y%���H%�ľ�>#s��Ȁˌ5�q ')rE��,%yB=X�����l��s���V�nH5�$�I<�W�������7�4�7g-�����x��k�qA���'�
��1��t�{0WC�x^��4'�~�k�R�y/H�z�'��P�g_�Z\�L�>0s#�w�p�9m��_u��� w�Z� Ȉ�S ���P�Uf
B��4��75X���H�*�3�tHi[���Z$��k�ugT�-m$"ܶ(��	��.�T�+���r����Դ�	a��hi�Z+��"�/�O��+���t�X�T��[��N��ѡP��]���1ŏ�]�� �Q�?Ɖ?Z�R��z�RP���CM�����LH�*»�^f	=�N��	O,yn��6o��&m�ub�F��ڷ9���ݒ-�P�h((.��Q��\��(;��#%E��	w�:X5�rv�� m���
5��S��<�<��j�������F�z&PͧK.A��#-q.�}��ͣ`ںx#Ш��'i5��Lf��t�n�(T�Q�˕`���09��c���Kg�������$~�u#��1P�7Q�C�\4Z{�t}v	��]P͎�3�d�M��[���0jzA�컀P�|8tmU����^�Ab�k'0[����O����	��z�q���mP��_V�A)^���Wi��w��X;[;_t8:hFB�@��$
��S�np",�`���C�}�֑�1��@�E�/#������fM�_�@�����7�g���HK�?]��yi�t�c��#�맚���,����}EJ��� �R�r7_j��]��83�
�HI5U�2 �znzs*ele!�=��+l���uL_���1�hS�U��
m5��u��%��Q���E����M��+�A�&��7.����(�.̸�=*܌h��:�m�������S ܎�-���Nsҡ�]�����fd��*��Ȱ���.���"�v8��n�hw�W�9��Br ��4�ٯ=�:8H!���wK�����.p������F�����%v���T����Y?JTq��9.*=|*׳鿊5�AR�M&���'���STxuE���t�9�\w�r�BXLl��D2����@�P�ݷ�z��.Z�]��D��O>���8��j ��_�q��)�RØ�|�ͥ�XV��'lT�+~'���T+cI�=�t~�'\��u��0����^��#s8u�U�E�<ȳ��~��l�T�%�����͛q���9T���< Œ3���K�a-av���,���m�*�ē�aG~W���S4��fzF� ���z�������Ԡ�E��Qd��v2͞�7*�/���q�	b�G�`��Rs�	,h�Y��S���2�Qv�x&C�B3v+h��9�����/�ǎNg� �WP�sk�?�G[fa�z��JX��\tW?���j�_�ng؞��'��iM6p<�E2����)zmgc���>i��N�M� �C��6`a���p�!�\^�Y��
h� n{�FZ���ζL=���nP�RR[F��^�T�yk�Ɓ���I>�{*Әރ�1� �x-��aPEr�J�7�c��o�J.B�����cK���7��A���`��o~)�{}�Ⱦ��{���[�еq�J
"_���5׊@�V��m�oD3��[4��C�-kR�
M�}�vh�#`)�`���1�W�� ��Wu�`�k�͟�i�~�}`2�*J��#&5���h�]��MY����&�Gh� ��G6u5B�O)O��'�Q�hX�#ǒxR�w!V�w���/���v_�1b���u�
�ܺO�F߯pQI��Y�ƥu7��W���B�D�Q�q	�qX��jS�\�M������r,󾦄��$W+�3J�N^4Q@�a�x��IB��C�C���I�a0+I||���Q���J7���dYĳ6�"Q��)�DU����oݹyb���5pq]q�U�\������H�XF��B�%P6Q9j�n*�j� �_r_�
%J�F���u�g#H}} ��b�I����j�������ڞ"O*V�%>,���u���څ�h���̠�Y�a�5\�DF�Y8$����hl[��O�eiM>���G��E���ė5����}kng
.�(=nAe7d[��8��$G^gR\x��M%��Ϝ�@�dy8��;�	�>���2�7=�K+���:O7�'�ﹺޠT*�W��B!+�zњ%���n������`p��������V��!�+�盂�HO�d	�QD���-.�ϣ�+��j�c�5d�yJ$���#��fk�����e�?!�U
�����Om�;���!��!j�F���*���q��/�P��M{Yx2R	�^�g�ĎMkk8��U�&�H-��uX����J�YYCa�GC����zq/�s7�J^�4� 3;�dN�(%���H6o���)��w2C��:M�޸d��zޝ�>��z���!��S��A��'Oq�jc:��݇�t�6!��k�E�"Q~ąik����cz�$�;�Ƽ�̪������̆��<�K��]�H鋳N%N;�ǐ}Z|A��|s���g����W1�S$JfV�y��e2��~ @���19h�����̑q����_ʐ&62���>��cf"pG��ֱ����ǄE��l������c����_��M���I*���P(Q�e���`�%�� �������d&���ٝů�wB'��m�j���TE�����.��Yl�x2	|���%뗱������,��{d~N_C?]�`|מ�`U~sU�;�=�e�P^Tw�}��c�m�{���)eY�|>p�΂\���9�B��DV$H�ϖ�.�5ܟU�}h}���H��M��б(�l��6ٔp��+�����]��r�b�ʭO��&ˎ��p�z�T����IR��/L�2B{�֯����`����y���k̋ʭ{�=k��b2����\�������o?w�5q�iv�0��8,$������U>�b�<<{J��fry	&O%Y��!B�Tr�3��Q��K�������		�lCT�m"��}��a��W%��f� 4����z�E�2��:¸�=�i�>��ڈ�{���b ��vabϳ�ߘ��+m��hY�N�+�P4_8l�N؁���o�(��TP���M��^(��:�É%IS̬Q��8�"{�v��OyGԇ�D��"������]��|������tvz���嬽�/��J�Z��4h�)*_�=�yGb�z�L�K~���SzyVJ+�������dJ�g��f����ߓ�K���9��$ yH1�v�';���ĺ���Sj�Ƽ�fM���+�����ZԀ�"��[+����"�5E1�p�m�^V���H��e��bg���Rq[8����#����]���Q�$�r�MZ�.0�7h�I�v�ԅ[�4F�P����`�� Tg�.�����J+�t!�B3�q���c�(����7����k������|�a|�kk����R5�[�˴:o��f�x��(K*w��8B'酘�i?�;Z~�<���'J� ��璫W!�lej� �4�L���L��಺�ߊu�/��$���9��(X�2��m�S��S0�	_�'`��^�vp���=�s�yM�t�k�C���<$D�hxd�$����U
)O����_�>t1,��r/��=��Z������ϋ����)Pؕ~���:1Q#=vH������F:��@`��W>�l g��=c�����Zi��Y�o
�X��6��<�:M�h���n�8�HLYgS @\���	&'�wa��'�S��H���R�9ƨ�5�8_&��Vv���[�I�D-o&u��Q�������s�h�R+Kچ�n�R��굕끑t/[�G�X��TZ�7zJ���L�BSh�D����$�c�C�Y�a���R_s:���yi��{��Y�g�ז���f�:R�G�n3�heP�v+zc�����W׵S����gw�CyUH�|�MG�Thઁ��3��Nļc5���Y讹LiZu؈N=5	5�n�}+�,���C
:4�יO���K٭�E���)�<�ES�m7��a�ϐ��.�>|gd�C�B}�,v�?���_��0�����$\`���|">�-p&��>���g5�C�WM�8��5�ć�Ʋ$��К�'��^O_׍�]� )�W�C��̈́�9����O�Z�!�q��\lV>1*:?�,�gX��GiK�JZp�ʨ�'��TY ˖��-�:E�F�އ]C�h#���3���A�Bk<���;T���S)�� �����y�S�`�&��{�a,���",Q��𤾋B�v>��}�8H�DR�AI�a�sYDXA�új�1��M��E�g4�RҪ8�n�D�+,����g�����q�����]�(k:�w��W���;q>pS�����(A�O��y��~����%�ep��s�YЎ _��uB��Ku,}���a�6Dƙ �[�+dw߷Wa�\볚�xp�L��"��o�~����v�"뱅Ɔ�I�g+�h���f lEMCK�
e���;�Y�o�M���YD���G������K%���>]��3��A��V�O��=���@�m��+ �ԁ�6�˚��	r�ɯb��c���t�/k�g�tǷ����h�$U���[���UY�U)����:钥��Z5!��U�o\y�x�\��܏9�7K?�����1�3�i�a����յ�y0b�"Ѿ�=9C`i�Ռِ{ư'���ZL���OR�?ԣ-�yP�زP�;��\_:�J��v��a\���Û|<��<(m�BA����$���VLמ�~�'�2�x~���R�X.�>��!������*Q0�(�m��S�o�>Ň��@�S*�dn�������}*n#�v(lq�5!Xp1��ʅUw�_Ss����=���,�$(��	>�z�qsʅ+ڒi�n?o���,�|����Fo8��cO���5�t�6���KG`|�CjC|��9y���<�)�G77+�y����SЙ�',��~M��j���,M[�HN��5^��Cs���2�������@X�|�d��4b��x�Y��k�W>�n[�.p���[k�Tbۣ�.$w�PX�}Wo@���cB��R>�lQ�ڒ�A��t�A0�w�˶�0�y�0��y�Y��3���-���u=g=� 	�-tS.���,�Y+Q�FX$OѢ��.�Z"� %X�$R&��2倬�D= �Hʰ�UQ�QXe����0I
��[��#��ʑ��L��
�����i@A�6����d��kt�O�=֓¹�.
2�T�'��Q!���N��nN���G���qw�'�w��ޖ�YL��q�ly���o�/Bs�~��˯5����*?%�y6���ۑK2.����$
��J�Xc�_��p8 ��m��8�����ӛ�5ŅͺXSQ�}_�Q��A��^���w�K'�-��d��6iѮ<�'����<f�ufToP��W��+��0�a;�	�?ϛ�����Ͻ4�
 K�UC�m�;4���R�@'Ï�MBAc!ۡG�˕|z�K\��}W��F&�Ϩv����w[���������'<��O\Y�G"g��32 i�K%�d(sKl&�@q<[�k�.�TN��pɱcD�МH����[����)@�!a��]dV�]�+ɽq�_<������J�.0R0�Q���7����(x�0�Mk�f�,��՗[�RD�h���F=��(�d�|=� a�o�r����l���$Ɛ�f����Bz���h�7���/ˡ>�I�&w�U��b���D�=�3��D@�����Ո����O�4z�=!2Q{;�a�$4(�IK6�����8���pW���&��P���h;a[��T)�Q��pE`����>_�1
:I�@�N��AQ��dnϺ�%��Ѹ�h0Wh�[#=/�Z1� �.� `8t3x`@���S�=�|&6:]��Q�J��[\j{B�Y��#w���#�c8�g�.b�H��܋���2c6�n70*^������X��|�ܕ[5�_(D�ϳ:I`�X2�\��)���0�k�5-�2-��Z��闑Li�J,�P�Y��}�4�?2�� ]��.�ֻ��Tހ��{$��ֳ�*�vw���!ݱg�ņ���������E��(�����g��7J�t�?���A��n��$�}�/�O0���#��0v�d�:��CH�a���+C&xʮ��~Ag�<���ʎ�X$�Y)�H��ru���?�"���[f�l���C�)�����4��S-yTeىk �c˦>��������e��T+�b݄�"ܯ��>��r ���.�������^�=	H+>�D��/�2�tUD�t"�o���|ۼ42p2�K�b6Pկ=���ޟ(LH�w����𫉔�-���)�.h�Ǿ�"����/	�����OB��ۿ��]�3:�c�����d���
n�q��������#c�&�~�u6z$&�sݹ�)�R�������XZ�%c�g�YWe[��=�\Ju�`͒�L��K�U���^^�>+���ݮ��Ce.Ƚ�,�]@ ���İkwj��41��<��`u?k��>�Xæ����m�- ��������}��]�A�!K�,U:�S�chP'��]S���Nܻ�+�l��gQ��g�B��;�hE��=}��"$Jߜ����E�2�b�1^k!�N�I!V(-�Y��s�j\߲1	[]NOŏ���<�E_ 'S9�������~��A?ч+\(���j �8�$�s�Ie�|?
3��>[�'<��I��vD���X
�H�4�������4m���ۘ/��Us~l��Ӗ���!�b`dl�1A�X:h�.��!�Xv} r�9�Ld������Zo�F�m�m��фhS�]��H�jY�@��:+�Z���+1;�����`K���H�7(����5�O)ː��h�\�l��$wb7�3\~����D!���Џ`=���ޕ'�gυ.A�����Z������o�LSv?2Q�"��x� ��r�L�0��gw�F�� �:�fMr�}:0cBDl#<F1�����p}#�DV0�қ�im�S� r�n��F��3�+�����es}q��s;�$���O���^8�1#2ɼ=,���cʀʜ�`W�־5Kzh��Ǆ7�/՛h��:�DAd��Dr����9Čվ�Q�k!8h�F�<B�&���c��.�[��®�a���Ev�m��ߝ3�тWw�Ő�iX�q��.���錄M/ܑ�D��A����@�$��W �����i��[DW�h�{�EZD������8����|	��sp��s%�C��k�_��s�B���Q�W7�<m �%2�)�}�i����{�A_K������8�����s��W��f&�͵��=-sI��|Rh'P���KZ���(�{;��
�V���]�@���_+q�S��(��U�w�ţ��r�jdi15��,^���e�H��(>B��k'�����Srq����*�4�{=�