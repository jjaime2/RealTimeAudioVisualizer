��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S����%J�b����j`)�u�B2z�l� ���#�p7L�7>J�ו4Ű~;�W�I�]�Ec|f�)s��˓ߑY�u�����|��
)��0fkh˔#�v��b�ɸ�* ���g'�����3�93�w'�%>~07�I�%�E�v�+J���q�[���s"k,B�ɀ(L`C��E��"�*KEBA��y��g���$�~mFy��X���x�,ᾷ71mѡ� �<:% ,I��nu�t`���Om-хb�:ǬۺJ�:��\j8\�(�_�Fq�֫8�+1o��3�p��]��ۄ�Ұ�"e�0����G
lX�y������ͷ�TQ�' z����y��rG�b�Wy����N�
b��W-ro��7yΓL�@8;6G@E;�9 ��d��$l��Q�*�HCP����$�
Ⱦ�d�P�F
�@hg��f��}�b�dA&5ݯޏ�	O�ae��2�m�18��*�R���hV��@�԰8"�-� I�δ��:/ˆ�5%��_ _ ]O���8㕈��\=��9�9�-�d(:�w������aH�L��e�T�/�W}���yZ���@d5��~�[j���I<6��p%CְN4Y�sβH�Z��KJo�p2my��ݶ���������Dm�J�
-�~���L49a��2~e/!h�zy�����TWy<|����M�o�kl6��nm�P
�
�U��1��N��<�4��������k-X����Ug�����-�Ņ��LB�����M�_sHv�#��e��Ygw�xh�ٴ��%�Q�)�uM���fi|ӣ�˻
��Ҋz�IG��Է\���`�݋{=���\��7Ţ���΄�.�~�Y'=�m�)��g0�'5b퀞#��֮�5�(%kR�F��	�H%e���A.�̂�`�M��!���p]������'�	�\�<���%vM04�_sIqg,ͪ"���7i�C����/�$�X�}��qICJ�r��o��Ȃ��=�4vK��I$�ek��ƛ�`r����{�*\u~it����oJ;���H8�u;�V�Di?����{��{�c-q������M��$�^?gl���L��B�v?�)���r�7W���RM�k�-֘�5���,ek-ݝ?1�������F��,*g�;�Gz-�x�v/��Ϣu�ZCa��+<z�zh�R`�tG��R�Gz�]B��ʐ�毠���1#��H�`��f�9�y��dy����{�٣�L���nBE�\�s?��.|���Jy]���n�^X�.�����Z�{(h��?�����>�;�j���n�I(�q���XD��_���<����vbU?c�:=�/.���J\]g�Б�+et���R������4u�u\*1$�\��8|k�e&�Sf�P����6fȧQ /�Z�.���{�.�S8�C�6��k����p�ʽ6�%S�R����?f�Tx�%���������u.�C��|j2���9?-����s��1AmI�����'����k�FйM���3��.O"�bǝy�5T�_Z�5����ؗ�F��Ϝ���Q��Fa�>�O�[-v���=c�iv��i�|o��DY�ER6F[��］@��4t�N����,�����
�ѯ�������>ƨ�(-�)�{��hH�$���>t< ���-�		��=)t�N�p���>;��JA�6SZ���ۯ/��/@���@e�S�,��pJz��|�`���i�U��Q\<T�՟�9���*+=gT!�aA~'>������c���/[}�!��`}�xc;���?��� !��i�M1q�/Vr���y��u�/���<�~��c�C�:@B �&?����43�naZX��c
t�$��h�9ⵃ#�q�}�����V⍮���Rٴ���4�x_+IVl���z}E��hn[fq2�b�x�s;.�'J
��Y]��I[��4�9�AԘ��A�(a=�E��(n��E߁ʐly�ǲ@de||䋂�>i�VE��"Y��pPӲZ��A�S �W�B�5F�����Q{@Q��s����A>G)y��{��Ջ&=�̊�XO�K������6J��]s�QcE#�����R�]���>�5�|��ڨ4j�Щ�O��o�����O`ʬ�{`1��Y07�Y�unW5y(���5M'�}���x-��WG�M��73�~��J�m��X��լ�v�kc�as&���Τ$����E��9��e]�neH'ϱ��Z��*�ԋt�W�0���8p*�x�\��n���B15���c_;�b�d���7b��Q���2,��^^��8�g.L}�u!4��(G�~ ���g	J�/�~e�m�-g�|���=Mmo�_��-��$_��^FI����(T{k$qC�-� ��\"�Y)��[�����l���v_Q�o���F�_�#@b�C$�\�ŷ �Z�j/�ͭ9��߳�9 �����E�*�	�:i˯@7w`�W��t6��\���<I�&�� (9��D���ؼ��O=p�� V�N�ʄdY۞�e)�u�,y. V��	U����	5�f)���1U���K% <�&��:,�n%����	���S.��o�/����3ҹ��̺��uL�yEgAsbP)�/\��#i(jdSx!7��͵1�������� Ή6U���0�?7h�d�x~3;��Mȕ��J9�+�/.�rB�`FE�)K��I"��i��R�$����Qc��\�A�\j�7�e������ڰy�����bݐ������A+�}C��dQ!H���f����̝1'�;��/Z������ƙ��Ǩ���y�^��=�=�W�*�G	I��)� S�#wD��:�(
�Z���<�*ʘNN{��=����ذ�n������j���������st�Ru�`�sP����H8�L��tk�G9|�m{�{���*�m�ʟ+y��;��b1�@�ym���'���A��⼖VUc)K�n�eR�{�*��e���su`���)16��D[�3��b��,����~�����PzCJK�P����67Ԉ��`�����E��}���B]�+��Ϙ���]�y�A���{�l���W������=\Kz@��dOE�� �����A���O����Z7�uw=Ģ%����7&�+����i����Rҋ��b9�0����b.�C���W.����)�ew����vD�~F�������ڡ�qP�Mr�����q_�%�%V�j�\(�&�c0!6e����\4{\�	�ӳ��5c��H�9)��͡�~)��L%������h��G����T��
VÜa`9���gc��x��_��0J%6a�Z�>瞶V!?˴�8�b�eX�)9�5�gT}� ]��r���<$���-�ﱔ*Jg5�O�M����'�Z�)�]�XY��;U�,r�ߙ�	�Ԇgd�7��i��&�2�A���7�����*%���r N�w�U�j��,aC
b���$L�]�J�
�aFa*���e�&��e��
��zovTH�����l�R"P�5��M/�+�1�H��� ��⼤�Jr��$G�sBa6%[�t�F�g4,�oӵ{Ru�ka��M��vB3G��A��Κ�u����a6!gt\��?�p�����?�pq���.ӊ�V{[����Co��=��3��P���%������"�:Mհa.�#������Fw���򹄩���խ*����4��I*�%܃��[@^>4�3�Y�jx�B�Gܢ
ϝ
x��8$Fp��D�?ފ%��8<_D��X����������?�a��R�'� �X/����T�m_ɘ�/�K�1/*��s�L�,4$��wX����.��'RY3��8��qsT�YR#$��R*]��I�P��5Fe�e1$l��2O�D_͂J�6؝af^fv����!	+7��\!K4�;o�!1�f�;K�������p?,�ycʷ�{I�\��ȈC����"�% �Y9�-��'��&����Spz>�ܮlɏ��¬���l��S)�cw��Xj�߹%�#��r��>����Sj��rY$�}K,y�����_.Z����>"a�<ǌ�V���5 �Q�}3�����>��S�N�ӳg�c�=@�����{�I�;��գ}�-���R�Q�'rX(X/�8�q5B@����܀ 5&oN3�D5���2���G"՗�d�)�zq��b�3,>�VB�8��\���k����3V~T�H��u�h�j�h�Lx ��nB���-"��)k��N4�=�=%��T��Qp�Q�Dj�]������"��S�i�Y�/h��`�u�5q⫟Hœ?��f|M��zcx�IL���TA�O��Ž�A�)����.��f�} P��u!��L�y��ܗ	�Ro�H���(\9��7�q�G�na�����<���H`�Y/�~�==�&�ֲe&aj� ��p���q���f#Ypz;ͥ/ǝ?�'9	�-kz���Y��Q�O�l�1k96`�^;ߚ����+Ϋ�6/��ҿ����+�'a;a�sr�cBE�{���<ƅ{����8_)n7�h���z��5v�����HŰ�;�Ƿz�-��7p�3���4�Ă���5� t����6�^����X���+�]$`T����^�	�Tը=�Y����~y �?jC���B.���G&A�]~�d��E\���N;�g1�c�C���i���Ӫ�#d`�cN
P� ��zߺ�u�*�/�/w.�~q����ke/�b*��[�3�:PI&�L�<^��B�-�����؄�T�}��i}3�5�Sa�kF^���v���d2d��*05��l
��$�Hz��=��q����{�/f��ó�W������ �Q�Rw����UU
�{�&Z��u.ӈF�ہ��Y��VuPC#��v^}����UM�s�  �����G��o�j���T���P.���*���9����B:�";�~�rHmJTX��-b�I��N�jB�Wp9tI/���������G��ym���w�?eH���1��8�и>���z� 1H�?$�/����nð���P�9��������Ap���QGŐ�����A�'0�(���0ٜ�#W�Y+ݒW��.��`��ÈSJ�W���M3����f�'����x�K��X��n�#ă��o����=����fG��,Y�mTs��I�RT��nfy�ÛS����M�YR�@����`���=��l.��,����Q� �/�4R�.K��!�~J��gfs��h%���<SL 9S�J��B{��4��|�mk�v b�)l�%z��E���xjU�{$c�+���x-��؀���,�}�ܩ����G�͙Ծ��d�S@l�N8�*�3{j	V¹�\UL4U��(8K��c�#�EOP&4C/�C�؞2��[�$2�"يD���dG�̕;T�w�M��x���'O%�����eoZ%&�\`�/��<O�;IL�F�Q�I6�B��Յ�#;Kg�.䫓q�7�8���jf��/"�pg��@t���Z=@<���������Ap�J���dLQј2wkŌ�JW�?O���(�`i+����e|x�R�N����%5F�3�D:��6U�(���_薐�J�Je�C������P��|_��Rۤ�Y�&л�S��8KU7&x[s�6���X��<��Ͻ��u�r$�AQV�c6�pt��'-rg�ױ�o��|l�ͅ�-,\��y�Fz��&���!1BM��ړf�S�?_��,���F����だ�*��F%)zE^*ś}��BoӠ>�'��ܸ��.l"����t���\���ڬ�*�tN�t�y!y��ڑ,R{���gd�>�W�Gºq�t��a���:�&��X�hY?�����t�����kh�����u·�en��%VR&#ѵLT�ހ�0hB�E�n�Hw֨#d[Ru�
��1�/_�e)�{,�s�}��,K�q�M�/|&U�R��v.o�}+�&aY����RQz~'@�v�쵐+�\?B�� A��?@�K粥�N����Ew�>M��L}�A��
�6~':-�Oq����5��A�ũ�h^�����gy��㞹|3��$J��6��Pk�I_y�}�/y�(��wB;7L��sg����Ĕ�#�q��Q �ש�nt&ճ�x�P��Cg}�锯/C�7\{ɧ���#"ˇ������������3�� ֤E���͆v=]9A��j�?��"t���RT��_1B]��P/+Ѫ=g jMz�&Q ���,��#&y���.��+�����z}}J�2rv��}��\���p۶���0��Np�v�Jdx�f_�Vbe@&w��>�7�<����w%y�~�KE���`�i������@%�1v����-D���{��k����'R�o/9b&��Rn�b�A����y��eƑ�8߽5�W%G$��7c@�S$yK��l?���\�2�NÏˈ4�p~`vO�Z0G��}�� �wn���	D%S5-�٨1yW��u�{���h�baq��R�&iSEh�]e��i�b��d��f7��^th�+�Nh�Ʋ����$���FQ+��Fl�/y� C����]Q޿���>h���W4�W 	[x�:S08Jи�6*����r!ll%�V�d��]V&�y����!��j�÷��`���A��{~碭0
է��-tI�q�b��1o~�g�_����MR�������Ze�E��)�[+!�@u���� �6m��x
�e�����k��_�'���o��+w�b�|�ևr]����*߈�id�r��m�ʘ��=����F9�Eb�B1-һ�
VT�f^�-���J|���bG��L�b��Ĉц\��I�a��������2.Y+��n�����(�ț������� z��C����2�)�~�֎�[jv��e�kiyf��%���\�5�f�C��&��a���vD�D!;��2?hC�=O���4
���e5�>�6I-�7�L�g�0��S"����_$傂����\�R��}�|�*L4��k��+�h�<����&$?�Q�q�6��!�����arȟ�a��p����rk2��b�1�n`���>ط�9�I��W�p>n`ǽ$q7 _�X��
�d�ΧV��rT�V���X�#ׂ�G���x�g)H�H��}oՁ(�{�v�e˽:č\���TX���_��"�&~�A�OH�1�ba'��w�z��t��g�9R����f�������[9�9��Ƌ������m���v^;�qT�(�����I�$h�\����-[FF�z�+߰}�v���1L�Y4�'|?z	z3~��yW��,�"�7�a����&��dst�]��5��w�(�Wd.	���Qm�,��0/l��*�4g��QC���k�*��+�$�dj�ȿ,��L]���貛�ĸe�aE=���T0��Lt���33�������w�6v�xǊ��C�g[(�\�	�`-��m�S\�?}�ڤu^:船i�n�;}��Sh:l��+�q�-�V�	�ݾ���8�FE��a�q����`�^C���~��+�KVb�Mi_���M2 m���ҚCB0�����b��d��G�W����n�1yi���삪)��!O�!�UaQ� ��3$-Qw�@��N>�/�M��Eag�Q;!��5�7�d/,�{�T� b���Ĭ����	y��,,����͛e�F���zG�[������v>��6@5�G�'�Ȟ;'�-4)+�
��o.�� ��N���ů��a�C�ZN�����M[�O�J�%�}5ݡ	ؿ��9	�v�����o��)�N����/��'��ר�E��R fk���B�͑/�d�?5���޼���Ȟ�cTyw��4ܶ�Il�\;#^~��(7�����.����kb���W��y,��3���#]�hs�E�d
iɤq�S,'�O�qD��mo�1�ԏ̶�2�6��E,��窾Ψ��T��cV�{��%@r֓s�+�vvw�R{���\�\爝��x�jr�+n�I!RO�>]��k3��4>�l��݊�Hү��Z+�3�K��3�.� @7�7���I������\�k�,'g�9�"~����ݐ^;G����ѽ��/�b�Lxȃ8���/`�:�n�R�)M���8�p5�Y���堿:<�K9�bo�$%іl8凫D���֠K�ETm�8#�3�����2�k�l<�k�:���.��N*��6��hj5E�]�����fnHͣ����AX�>8$���wgk�ba��9oD�!���Ǉ�md�1��|��?��BQ�}��{���bLn*$�����P�a�R�z�H��82"�2c=�'e��U!l-�Gej��_�-���t���T��|��
|���pa�U-�i�߽��X9��o����@���}�sO�eZ�V!�=�d���.�T�wrԖQՅ|f����(�k���]Ëx�HN�:�9;QQ�����!(�o�����N�@(�m��iq0�Z��އ�r� ���F�*ڈ���U�&�N��q	��������P?�~��fPD�4������v)����Fm�u>Q�<�L�D!��],י�m4��,��'����o(ڳbU�Mo�H�����p*P�1�F���TS�.�2#���A�w��6��3ɯl�:-r*~�q,�����׭�Q����|�;�h�;?������&Ԃ��c#iO_�^	���B�r�2nus}��'Ѻ��8�!a��D�Y�[IN^E��J���ٕ/��&-K$}07�5�>��]��@pyX5��} �^-����{�9	Drw$<��34zZ�AP9���u�,�b��qփ��I�:)�E��M}��Uteڌ����h\%s�G{ѕ�ed�裧Vˣ��~�6ǂb�b rY��[r�x'�.Q�9�\�҇����̊�J7^�"�|�^)�����4F�����b�##����m�Us�K��Sb�-3��0(�d#9j�0�>�%��u��҈�t�;{�o1�Ne�]��nn �_��=6��p���F���G���^d��$�Qzmґ����t�&�Fk��}|1��8)X"N.qA,r�KP�1��f�D��>W�'�������v�2�e9`�eʮ�ϭ�����������y��F���M��&�H�Yb�M�Dm<bmT[�*�(j�d�v�b����Ǆ��s��"�3(9�{
��ci ���:�ca(��������:h���>�gٙ�BιQ��ig�.�K�Jp�k#���:F����g��0%K�R�Q�.�����{p�Q���-K̯�ń�K>ַ%È���Qo�W��]7�v�ƞ��Ox��)�VS-�\R��V��H�R�<��G�+#�@uu���yIT���c������S�K }�$�)�����JA7��4ޓ�.�A�q4��4}/y�o���I~�E��~��xcr������a�"VԈl}�]`�������M�mR�� �%�=UH_\A�80�*�����p;�U ����v��f�0�L5$꺭#=Ooc�:�"Dx��}����L�}����uΤ����N���ȕ餝0׬c�E�'���U�����˽7g>��`��� ?.�,�o��-aPz�!�vu�����n��W/��˝�?�?"Qoa��i��b[7]k=��Us��а9/a��ڝ�eF�&��3t��g@�D�ƍ>�4A-�Q�uF�Տ�y��p�ȵ�;HTaD��5g.���⮊��j���H����Y�=cg�M� YSA2G��=�����-~��G�V�#s}�� 4|�d7���%��-R��1�w�i��/��}#=H�2q�v�/xZŕ�U��mm��`��:�U�T7�و�e���E�%�:��2��@���'}��Fh�qu�P�FOW�gf�$��
�����p�9�$ى�Y�!*�<�_�����&�{�%��00��q��xd��L�ڔ2�к&IN���$�|@��0�~1m=AY[�v@��>�/c�ðO}ɶ�}X{���=��4$���-�J�xa�"0�~]�Y�D�|h�5�M��r��7Z,�!X}!9��Fp� �y�i���v�v�c�ao�˳li��%?U��F5�;���X�7���X�k� �s���E������T:B�	{�Q^���a�o���1�ѯ��������܈�z�X��vP���#/d�:~����O�嶀~Cj��J!��w���@hVJ��Qq�{�U���CDJ��J��j~��+���N�t�VXmw-FCa�\�@�<�˙94�ώ�0r���E�G&6��@_�¨(����r�:��Y,`y�ґ�ʝ3�r��p|Q��Q w�'S�w��,��&׸\�]q��8�&.�?��V�>.ͰLhݎi���dᛉ���>7�F&����2����f���� ��D�����U��)>�E�v�b�O��%r��z5X�fڛ���Na���#�,�9�k;�u�26y}�^�
�!,���uyܮGa��<��wSQ޳��2Zڍk�SR��L���Ul���d.xq�k��WCl�]�U�4��H�NOXK2�B�4ѨY����a	r#����L����\�	!�v����X�W���s{jL�^�����e�9�f��o��t-2�80�]�U�l@ӹ�����;��xh��k��B�5>Q����x��ɼ!8��*7XM��i��xu���A��)��LyR�Sf�i̿�
q��UM��\�A@iЅ��<�i���:�}'�>	~���~�*	�)>��f�漈W�]*���W�����`�Du�s�s��c�k�7�}�'��w:�sۼ�[�&�� ��V���s]/�4w��s��
ı
�.U�!ꐵ�⡆%7�@u�M�4R�bv�9��q��FpY��a�1V��8�D�T�E�<�	��K���T,��N�y2�3[�x�&��k�b�ȶkO9���A%��y߷^w����o�BfD�,�׌�gИ���զ�,���
Mu��U!&)ؒ>��T&b�$�k�^�b�q �zi5���g̉K+�n6�p򷮕��
>V���3�4uN��'Ѡ|�ٍX!Q��B�7���C��I��� K4E����wK����d2_F��ም~���M�m|���r�jX+ԗ9��G��/OlAyoKe� L���s���%���ɩTI��
{KI��c�L�z0zZ��8I߁�&�d-������.��%u7���6�$��#�ׁ9�<2��
! 5#�uj^�;�c&�2ƺ���*kl��*������H���; ���0A�aڡۚ�	���.�1�x�A�s�b��?,���(Dt�?Σ���=e<D�U�w�'�:U�{r��('�0A��	��L6�F >�`�h�'<�I(�դ�_밫����;l����4Xt��2~_$�,0����G����8��.�v謿	���^�%�To�@'ϱ#��y^�G٭;Erq�����C�^8Ѿ3I�Hr;�}��~u�Bk.��*���b�,����}o�uu^}���)��g�l����ĚGG�Y�*��
̚��KAZ�?�J�Ұ9�<�%̝��~�޸�^�Z���G-s��y��L� �SC�=o_�d��8,# �8�� Ӹ
��30v�g>i�6�'Z��W ��.�;:���� O��Yhyg۩�<�pX��vȮ9z'�r#&L�Ua+Q�J�u���F�}�^a�Id��	�d5gh�v@G�c�z� �ͭ�At�u����}����"� ��ݟ6?.+�T	�J��y-�	���U_�����m�u�Bk�>
/4���2�<IR���ŗ�Mk�A*�D/�#�z�j=���L��\ �5Q>?�����~#4�_��8R)*�0��H�2���ڷߣ��L�wS�L��l.k��U3�%�l���kU���Gs�N�����8�ͥ�yv:ؗ�6�t�G��+�+��P���j����&E�̫�V
o�R`��P̱�q����:�|�3q2�"!H��u�_�$��w>{&q��Y{���aN`�?�(�f��Ĕ<�����i�1�O.t��p{�G��J��2��.)�H<(߃����PNK��~��3��Bۛ�:��N1�#{�;D7/�����e��M�\΋�-��A$���P�v�0�{*�}�s�����^�t����$���Z�ց�G=Hk��I��S	�\2!���`��|r� q':&�B�����c�'���_՝�e���J%���7�p,
�%���+��Ж���59�
��_��T��'�����oґS2�Y�A�(�uC|R0ҽ� ���=�e4i&8�K���ў�i�������]�^��j�W��}��c���<��#%|H�����u1�d����*��Z�O=����:Z	��{{yX#�^�P��
�{Vxć�@�n^���r�H���E���c,�s��H~�U���&��Й�y���m�Į�&�������U�i��b"h_��x�����WA#�|��
I�7���"z�Cy�`*�Up!��kl�w��+��@�.�O�i����M�b̳KB���ZV����7�p1����@�֛ME鐵��м��*;Cl��M
���