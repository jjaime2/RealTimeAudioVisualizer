��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��33�z_�`�f����EW^7"q5���K��Ҋ���CU��ˑ�v~,�ynfP\��j��I�qS���=r+%T�U�o��I�y&/�T��W�O�2�RqmTf1
r]âN�.��&)�M������`��#�<ⷝA�.�O҇��{�hm%�~w�½D��t��kC-���_Uy%b�X�K���x�7�!+*r���tkO��0�[��F�B�ؽ� �$��2A�����'r:�8ƿ��fi[��l�OI@�� �H.��������}�BG�)W��6ٯ\��*i�J��nv��ٖ��;|�2�H�E ������,���� �+��ߦ���� TV�y�V��u��=`=6����ނ$��C�����m_O���׌�U��H�;�!�S/�Ec�O\+묤ć>�.uk�
�P��?�1ɱ�5h9D?�3eAϱK�����m`\�XOM*�����6��$�S���Q�p_sQ�";�'��6�i�p�LN%�*�����/��;�)\(5y�&����{����>�Q"�5�<@d��
�N�(4͈M2����Ĵ�*�8�rSQ�!-ՙ:2��V��Ϩ��@Ǣ�(X�M!i	-T���1�!�U�ٕ6�qL�z��8��o�r���'vi�<�1�B�w6���V��R��`� �/�8�I��/c��RD�*9�e?���ԇ)��!�$!����ۊU[q���g�|�"� ��n���pmi�����>�����	�WRȩu/і�|m�<��YRS�HcH�D���d�\c��!	��]�0@j|V�Pr�t��!�Đ\���ko�	��?"����Cg5X�D��W#��|6&���	h^�� �������vh&z�jY�*;�X�6�z�ց*Iវ�����9K�2�C�E����5��q�_���8l��Ρ�l�Jl�Jog��_�0����n��|�+>m�C
/qZiJ.L�ˇ[��VY@֬\xR�!f�9�0W� �āC���4�hqF٢S�ù�/,���.����������c�f�10��j�\O��+�q�=�mO_OV�.��1 �R�Ғ+���G�\"���+}dܸ�k�m�g�d�V̕�BU�
��d��hb醶eۃ����y��ah���1A�����w��f�/<,Z2D
8�`�R����5�n'VR����͕d�,4�b�L��0�9ߎ��}>������G�!��w�һ�b�b����5�˦J����4z�E��Y6}s�
�7�l@4p�����+���e}�h���t�u۫`td��aS��M�ȯ�������50	wz�D�p3��.p�B�WȩU�fx/����@D���MÈ���-�J�_a�M������.EMT8Tu������<��B���A`�}c8�dy����o甀3�}�'�,̻`ޝm�X$s�Ť6]$.��w@��b��>NW`���S��t��;�q�Sc�_�B '��Z�Q���&܊IY#Á1m$��V�A, `Ǔj"�x�xv����N�N�!�3,~_�+�"�Q}M�ft�>g=��N���q,|�<�13'�p^r�v�?t/jS|!'���H�	��s��Vyư��M�{�zN�P+�&r�t�,���e`��R6_�r8�KFnD�n[V](�eBĒ��=�F�-�������E�	�t¨�B���n5�?�;��n�<|�sց�nq�#���lh��t�����w��;#\3�8�{����g7����iF�;�Xф`����i��p~�3z��Z���3 ��C%#ĉ;�zA�f�ci�{��6�����C^���P����Q�T8��ՍqvoKb.V�⛌�ƶ,Y|x	H^�P�����p�Q�����|��l�=2^Bl@j!����]���v6�M?}��S�ENW�B�wĊ���}~*�ɿ��Id�m6~�r�0lEfSEsEO�E�4\��A������Ba�Ī�`>�6!�	?�T�@�A�ˣ�tw���_�2��Q�an�ߓ��
�)�m�ϸ��`��N���
�870s�z7����E���k���*��31�����z�~ڄ9���:�®q$B�~
ΙA5O&�;U��~ٓnq!5-��'�<�ō������}_��&���ش.�����&ס��=��):~���|�O�o��Ť0U����d�Ǳ8�X;�J,���d����9��u�_/pt�h���`NDJP�w�#d��֊��hot|�sp�<m]��Qg�~��w�K�tt�	lR�5#k<2C�P/T�2���Ⱦ�q���]�I�䛯"��.x��m���W���;�W&�c�����E�s���9f�kF��-%����T:Ҝ����.�����@��fxs�TR7�7>-܃�&8V�_��[ɚ^��P8j�sۚ�u���"��d�5޿�1_��d�٦�0D
��M����I!�C�*"+.�N�g0B� ���g�0��j�|�gH-8A�@_>�o�#�}%��)�^�W�M�;�Y�� �7��������+碨w3�۳��Et J#��΍!{wSBNvw�5�Jzjۇ�7�ƭ_���(�/Cm����x�������9�D�)taQ��8�u�b�Ԓ)+?���qFU3��85��GO�.�A�Wiw�Qq�491Tf{|Үp_�q%R��	H����5��n�����댐���q�4���Zk��� S��x�5��&ag��Þ(��x���2
�4	�7Y=о�`E�ڝ)�FD�WU�����P@��\�LlZ�w��:���Ӯ�W&]M���6�f1�f4@�oϷ_m�A����9��qe0���V��Jh^D�����Qz�C�4͵�)L	� +�d�-}p
0#֐�������т�����|���:\�x�S�֑��L�t�Rr��QOo[W�`~�X��ŸOZ��f�=��W�=3e�WNr���z��!�M^Y<�ea�t8p�1A���ƽ
o ?�c��5�eS�m�db�s)���W�e]�x��G��<w`ᠥ�$L��S��	Ͷ�Z�Y�[?��=.����e�/W_��!Z�A��wFg��ja�>�LR~h�p�"y`p&�ߑSv��3tN�e}	)h�"�ڏ�Ę\=�)�p,,�L�U�Ȁ[mQ�)�@�a�Y��(фif����xa��6�X{x��2�l�P:��V�q�F@c Ѳ8x��U*�WU�&L���9vNC0�s����y����8<fx`*��K{+\m���<�P|�@�y�'�,iD�.�!�o�L9v'���]�	b�Jo9û�3��ѣy�!=��}Q����`�)[������ፓ��� Fh쪬�Un��?`*zE��f3H����`a=?a��w��b�X���>��vj30&ՙ�E��}E�)�:BNV�@�L<���ܴ�X�=.�p�w��_�&V+I��r���(�xF�V���j �&�(���VcXVl��r��.w�gZul-�x��$����\�^���(	v!bU���f�\8\4��Mz>��d�|u��W^f�M��ˈ�S��{���\�F��f� �O.M���:�W��N��?�\��/5���K�օ�;G�!�R��Pō�*ţ1�Y�<�o�A��m���"*>�D[��_���`$�;5�J���&�c���'Ӽ[���J(��beo�է��A�ze��>��	c��(le����$���W��2k苭,S����h�.�-n�p��=����{���<��e0�Ml�(ݝ�w;&�37�jZ�jb���/�����@up�j��8`��.W�V������#)d�6,VJ�߀����߲�d�y�GU�MI�o��ӣ ���W�G��H�7�z/q�mr��$J�n�)ٲ
�A��qP���rϡ�`�5A^�
�����`-!��&q��u�xm	"Tc���?����X�*t��w��ä�y�X��!��Y��5��|���ۇ����3�Y��ښ�~io�&4y�S��I��g�c �F��v�ֶH�%&Iˡ�-U*��sb�w���]�B>�	���>�����Ŷhq��'�F�]�t���y�\](�E�Ȉ��b��y�\=�~�;y�!����:ik�2��������w�����O�j�9�	y,N�/
	�j��cb�I��naB��@��DA���#p���::�Ä};�$�H�i9��:�����*"*�(1W_�hǣ���`)5 uN�:NY7"�$�V�}����0��H8�~����;�؅t�&HH���%Y-�X��f�9�YVh�@����rCo)�WLD̮�8vW���3h@5I<T�ŕK����W1��\��\ٍ�VrC��;��.�-�F�z����E�����F�]�n�?���d�Mꈈ�G#A��i�|c��r�
�Rڴm�IR��i�	��r��IG_/�"j��&�������OWjGo�|.���a�m�/8�#�+ �%�X��Un�	q�E�����A
57�d�[��к��ݍ��WO�c�[����ܞ�1j�m�[
��ϣV8���|�ʲ�ތ|/V�}��h@�īPZ���9t�D[n\�4���`�<��Fm�tk^ T���	�Ƞ�}µ�yUʙ�p�a�O�t�Ì��n��%�Pm�!a �d��DWF��b�@"ӵ��
���-�`����g�&�՚hke�a
"�y������I^)h:Y�����&�ϵlrS�gό���TD��<�<TO�PW�fJE���VW�?'���4G�������&"!�E�I��w��v�02t0�Q�������|�.��>���'κ#��;ʇ I\ux�Y�w�N�/y2hXt���Ë��L�Q)ry	%��5�ݾO*(���%ޮԆeSi�y1-k����MΌԅ�O��齼�`��a�+y��R�u��;|590��.	���������.q��i-����ڬ��%
2�4����1�y��h��f�L4����������_<R�����T�@�<Йk�f�	�&+S(�����,_I,i$�}r��\C	�D`zB|w����2 [CX:��/�,�����%����S�������S�Jݾ��=�,������^�#x�Ks�����RK?�Uo02�x�L](5(��9�*u�e(�Wg��dȣ3M�O0&xvSu��q
dW��Ꙝ��]�)�퀢e]��m�;�C �R�#;I ���bD�c����ar��_Oru�Փ(��%/ gK��w�^z�4L��fKp�54z_ė#��\��$��;�UU6A4|�$r��G �<���uάU���Z�贞A_I���x�έ���/cy�UPs(���z�A�Ễ�U���e�����(�_6��fvpf��/?Z�=��F�K+�-����"vf�>5t�Z5\m����V�繠@��xu`����꫹^��{J���=ʦ�9� ŭ?��+�4F7ȃ�d�U�,�����t�#L����z��!��1�m:����뇧�3^4�2m|v���f�-j�w:x��-����_<]�рЍ��ֲHK��U�]�y������ b���Q����5��C�Z��Tz�(�Ђ�F�;�F	��
&Y���!j�5��+/+*���͐}<-�ɇ��Y�ӛ)
{xW�()֔��9��P�m���q"T�89
�Y��<�1�T��r)�Qc���;Ϲ?GY�G����Ez?���
�?�!��o�tpf����/��xX��@����N��������5���.|��6��N}1=�t�\�ج�ҕ��s�{&_m{^�_H��s����JHL#���)9=S�2E)uB�Z�@q��� ��G���\/$2c��+#D]��"�G��C���i�8�;*�7�{���*����z5�{�����E���AL"�,�4�>��Hٱ�n�|��3�뵜TsaU]�<���ZmO������3h�w�������s29"�Qk�,��3�f������ *��Ȅ�(_R`|����:�?��妯�mH_�mǘ�Jׂ�
1R���K���6�~:$��l���n�1'���`�r�Ӂ�.ڻ��Ĵc��d�9�Ș�����e���xr�(�ݼw� 0�R[)fQ=���۰u�i�͌�_6ﲖ�AwS6f��{�F;5���Y���U.���Y\�2��p��V�"
l�Gǥ�F�$D����T����@
��^#}�� �b����:>�i}��!}�\���e����ѽT̻�sy(а�Z�M�̮h���g)�����Ha��DF��(�4�b���W���!� �T��q�1��,9���D{F���E�EÝqnD�~�r�}�6�0H"׍���R��������uc��.^~p�w����j%@�K�v7�����5��Ò����*)OuL=i�x	�l�7,n�x.�E�0�t��?_�����-�;a���m ��)�$�Թ�m�Q���)5� ި�F��K���?⤯*B�_����i�u�0W}�IMDY��b�\�N��B����φċ�YL��d ���DZ}���EXj}#����e�\��+C��SO7qf��C�C�Z���,�^�I����I�d�C�G���5vP��P�!��j/
j��5����j6��y���>�Ӥ����⿒\�����8Wڑ�kJ�Č4�l��`0mã�ׯ���i4"��X��Ks�vs�p����j�x��}�����5�����81j(�V�")����YR@*|H�9���eH=W� �g</���DM�L#.Ė��Tg�^f���׵��ȴ]���/��(��̟��H��acEfC�څi.	�I�b���}-�p�;�h���B�%�9�=�����l��+[``iI�k"�y���ɏ��u�d=����g����%1�U�#�����~�t���b�m8��L�xzAM�c���or����jCc}f��RRy�- �Ʒ�+�m>X,�MT��Sqǒ���G�����)����ڔ�;*%-FHҚ|���0�M���;��}��f�T;�%����်��j���hOb�x^I���M���շ���5���̘�ǖ�G˭�c���d�5&UV�n�zm�<�h�f�I뫻�;0-�HH��0�q�U� ��H̀�wCt�̲�F+.�F[c������Ȇ�H���wqce,P@�B��Ic8uI$ڋ������\o��./�� ���@���n9��^�amV���7�pO�@�kc�F-,q����Q��V�]�l�g= �Kf�h�O� /{~�$�<*�r ��B݂E<6��Yk��y��NYI�*/���2A���t�x�rߡelE`q�W5�JQ���cQ
�����X����N���m!w'�VVw4Ql�����Z+M��*pQ+b��6�&��BĎྶ�M]Y��*i�����x�b<�������Y���ݭ���˹�g˒��0VزW�B/PHu[|�:��h~����R	��o�Ig3�o��(�ڝ�n��mH��%�;�в!���W���^nT��VF�ه�X�i��p	"�����l�ޭ� �-���0�&�F噿�"�ؐ�3�1
������p\�g��Q�p��v��Vȍ�2=����]%��X��֛ݍ����q���b������(�:��^3J�)	ܸ�6��15U_�?����A���0d٥�6i2�>.�PyHm�,V�́�$�L3��L�N�0r-�@xl,n�x<3���ޅ$��wJ+�\�J^�z [�$�j=ct��;��Im�NS���)�S}�<aKd�)���vc����Y}9� �J��cܹF���Ĭ_�i���p���h���0%�U��h�L@����c49�KWC��] �������됗�P�nZ�.���a���� �z;�����H���Jlַ^��bQx%�����k��!#�& ;�di�j��\��_���6iFnYDo�-���s�˜�,$]�±V3ͨZSOD�GC�f�1ϱ
���
;���hI�.*Tty�Ȳ
G�$l��,V�܈z����ӛMz�s>�z����:C��%�:�DX)@'�PK{A��xO�?87ZBBCAam���&"?ѓ����Oὅ%��[�aS/�3$��#��]�U��O�F��xN�8���/�fK8���V�wS�c1�]�;���O�V���>T�,Q�S/��}�}؈XLˁ#�7�F�(�^����^��q��(��{F|��D�?�RDV�@,m% ~�Z�Or�Eui7�U��m�[�6