-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
W5oYc53mFBNTgZUjB7k/Ikyws2R5M6qTgrxxIGjOtehIW15DW77Cj1WMpREFUadxcU4QcLIFErlu
+XYfWrOxR/T7dCWDwEEBLTmV1temdF1yk8kvEuRctdebqQtGprFz6VyOmo6weTWSaSCqljhmN8mH
sdlriDPfDz2eaUJi63DiaMfRAo+cUrzcxdF9H/A3oXFGCJ7EB9dsPOdiK7LRooErYIMvlmtkiv4B
ES9Des61pPoKSBNKxbM9J31ywpTtYzqXP7KFtQYhikk0yzaRO+hn+FsLJfyEstS+OEBGJn4VPMY5
1eiFLP+2JHY7UDaYCcKBVaFE16YNMuEt6vfiAg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5648)
`protect data_block
n+OyzDQfPFWllH6muikawBBCf1bLyWoMXdtcjLZqqF9dnTSe2ehAPgDF0WdovTtmQbpRxX/usSwU
sUG/zTmx0YXcNMG4Z2KTEecU82ucbzxZyVJI2Vg9yjpubaVk93IPwknXvJoJl4JJtXe2ShPnsbvK
zEaDsepek7YXaFxvZzfOlFb9VX52fEJAf8omMXOuL/QIiRhK1Sc5FBKK8duQ/as7Oo2Y0N6MwYcZ
Tr+y0KWghpqbx8F4Qav1TGng2pbIKhIBQHnBQuHLa1c2xCfF28O/+UaCi2MkI/ES2sxDUMe+scWW
4mn9cFUR/fxPnmF2DtJupf59dFNpnOmT3zm7rHj8tkQuFZsulz1ad9Do+EvZCTWjQdHBAr96uGB/
2moERlFtdrMDqqTjTwurs7eeEWn3NJxo8Uec8mHuagXam6l/ok5B1c0NYGrzsbxLDSiEhUN0N43Y
ukvc0dGLYC3T7c4zZu5uiJm7faeOHLxC8y0bhZvLIOwJa9SGdCiUwnbj3Lk96hGVaaDWlmb328b8
aVYwGhxlPLJzAYoTo5iCJI5nF39ROzy37p0wENh3ke1yPP+veY7qaHqE2sqnDuUdxjSeKAqZweta
1j/mrdjZ1Q6vg/AKIox5nGikcNs/PrufQb1WoVttJ/z1X5XB91rLevb6pvhO/0Ud6ClbuhndBaot
peQErfYEnMiA3MVL6/IfkcH9YfoDr+5v14whXmzGiWmbcqDBBFLLPSkN4ABN6EH4v5yuXO3wyHmM
W+VqkEMx6FgnL/2mfSP/ytQ8k3VqT+8F75vm3ADpiVZqztv5ft7x7x+LcRd/qghe31WF4AfvbYb4
eoHRfvSbn5ccR+xTLQw44ZiHhPj1H4OTX7HUc/CbphM81ESeeJRZcBZnJxQi2Nh0rCsQW9h68+Qi
NaXzh7TnQW7eDQ2StKWzd29E57gak0FG7Azfd1HWZeULbbctSx0WrLK9hyqZsRza41pKsLOZq82k
0HuYPPMNvPkfVbqC5IlHAFa8KYZNLxR3kg/VsfLLSnpZvtcj1DOaMCKSKa9qeNOcmmk3G/kKrBu6
KJt2wEWEQByfEBq1A7NahN2WdySA/m+T6WgTY7cxiy29svk9UDIa3Z1QH04dyeq2bGq5btS9nG8s
6doHap13/VUL/faHc/952+B/b9yIyBdlP8vmkroK+m1tNQm4XRXBxWxmeGAEZaLZ7VghUrAZkYcW
xnnJ0DS6w2QJRWyE6bU1SwmnDEVDRDECp+MvZclyXAXeWDhNc3CfLUA1pzqCFSQ1Lhrw75u5tYad
j2iwTi9TphTiY3WrmEX44Afmpp3xC8qsbWo8M3pRZKZb0FiM2LS8ylB/cpsA8dvU9oFeuty8DbDT
URzLchXd4PQpjxQupCMSeIuHtUeoBk2feQc6A7O1V0jlzqQOjNeUcvVI5yVhFDt8fXLMMG3tMwOl
hWAwBgE4hJekcWRS93kiJ5qWVK4YurqSDLtVlu2C184er7zgoG+xjv84SPBzZR9RfN4fwSx7eyY4
iFSJTdp9AlqFuP1fvZ7aItH8ARJbbNaTsY6q1XH+X0Zmi9z7ws/kLIIUxC+Pg+Qr1Wbu7xpyrwu7
S5ert0/uvUpvQW0ez+lwi26FHBD82MVlJtTmnIwl7hI6dX15M8tOp0o0EO3l46CghDKlWzhIwL2D
UG+o5KM1y494Y+dKkkx76LrqYSF2vUjA0kl6o1MKCH1OYijZe/qYTGHs+UcHo0iIH/HSpXGtS6gb
C8IAX//QnXBN0GaT9uc9hTS08WGU0e3Q1cIZDnKQzSvUiLCHrkz25eQ1Q0KScBiV61l1icUI3xMj
lbldIahqOXzCwPm6OSDwXBtCLYZRmHFcCmRmBbKwNyOEDkobJUKKHdsDEn99WLjsUu+Oxo4SfkS+
j4tB4UdTI2FqxjJvZbbgLHjC362z3Tw+qifWDUSs9CvAxfg6y6e5H/dNuUABFDE/ANVKMeLRH2q3
U+O0NTYfEOGz379g6je0SczCmnsX2lcSRLFZLzysQpztFhaNsTtJUUGGLho/i4LhFL7KNbEyfH+4
OkdkWxpYS84iDFXGZKXk1zW/Y1bN8P8HVAbj2YZsXv9mqnkHrX/yzszk2y7IDaUhKWMJI1cPnPEk
dU28XU71ZG4SEOG7h1GkOJZRQ8NzJWnbBDMDxjW6MieEoVXhXnD0hiRTs8MjC5eyCw6mcoUdV6pG
2D2rmkOQqTlScjwem+Iy4uipy1u23O919rMs37X2DIj+Dd7feDKYmIUtoRXNM7ZFKpUrN3tlWZ1t
vwFGzTCmwfe0cAPvXxdO7KrTVQYf+d3rn2AM9Ujpow5CQUgq2VVLxAA3YZAxVFV27OF9XWGhpepQ
eHSrxoIZkZGPOMQDHuRM76gmvbmbzNh7qea7tzhO5ZziqgjG2GaCxfgFh4VdUNTq7NSyw1z+NjwU
97JDMBW4IRs++GfINuKmUZIL2QfMt6MPm4MOmideP3JMaVGCjNpYAnz/fJIYE/oaAIWAc17P/tc4
6I2JZBu5Ht9LLrC4yzyqLjG0NraNZ03rbzRf57unWGnCy1CKOUrUuL0YpTLfJ5PZuEtU+7CQ+I1j
eOOgW6qgRvzJ+X+tlDlzjboIAPFrURkRrlr76OghWwp+lUmo+iYxGUxuzZu98WrgoygauG5oLVGh
pN26M2LVSEamlU7J8M3ZWoJ1KOvRWNDYc36uhBObrA2YRvIH3Ar47j6uaWhxgUBUc+218jjwDUWJ
sM2cYND/PoO1Klm1JM+9q62vfdV1SIjCMZxhatqIRwHPxH2OZ91SWLHcSRE0i2KTGaqNHgLPjAfH
UhLZsnA0UpQ+hQBapuoXANF1uP4QbpSdykYlBWYpliQuzsFGv0OrXplGU9i0G+7RE3IcyLvYtKZB
pyvOD9yLyxSo+tQjeMXemHMj8O2MuvFl/6uHRJO06V0/1L8/Nzkx0U3pRj1dTw+jH6x6U9iA/Kgk
rJZKZQVYbZtSVHGULyeQ7fKjH4NvMVJoyIOHwXTZIOi4IIByn9gPa/ctMW24l66oBfqv1rIlAVMt
yM6IwVmHAkFAx81PtQBdxvrnrgF5NaWHXZd+0va8MRh+rO5H/BlrT+Ij6XZ0seUfGaWleASZ900u
HzV5DjFGznL7oAN33BfcQJ70qN5Nd7bFnuyHw5+via48cJX6dOG6AEAC/LAJ8mDB+IYSnPuSaOTm
W59TByIDuYEWXCrZIqhMDn+VEs7KFhFYDDpW8usYGJ4XgRUY5XZ9Eqf66Jf9x6ffjFVVDdQlG3Ip
zjYMBK6X3eSNXlsh+fO/ucpQ07pVAMv8O/T0p4HSc2NQ3Qh8bRcAqNqWB7mL1NElKcq0Vq0Aa60N
EPtOXdNAljSuxmrx5ARSxflL3pDDjPCdsHDAi3e2fDNIyZMt9b/qXIIi4MLycNsjyuhV4pxUXoUG
xcGrbkjWE/GHnX7JBBRRIj4z+SoG+hBXC3p+DM5nMoRiTczuh271dexOQUmNcv9lcMRwpw00HAc1
ILKwvlvXuR9zE/G4fR+1Jt7B+a8frIVLLV7lYaGG7fO5E3NGQfQPTeIlZBq7yBUZHLmISAXXBn2W
GlqHyTJ5u6uLL1ek1FZpv+afFj+RW7t93/QOGjThyvuAdG8IIHJWmDbNX61a/YvRZULc4sVdGc0v
6sAb5m32vtHOSPbyS7o2oqhI5Ab6q2f/yKW4bVLY5/e0DoMXVu4zEpMbHJ9ATm+EbjuGh/gFjTBU
Vn1bNeCRhXPeQR5eV47zdEHKJiGUHj3kx5+gd1N+YMelzxeRH6QghdXrjeDy2je/JV1So27bhkrn
S/1Qr43FVUx+jZXT+dpWZnIOkBhINbtjCta8Ku6009GSC53L/dW4neP2539kLkQbV9rG83yKGlmt
bDwnDplQXqrt5sNl9qTUZz2i9nifK7S1b4n2x+bsMX6pesCBnp/+aR9fzSMeRDQAdhJHUgtOl8ZJ
LBSFcttQVHKCCn2lE4QGHXmo7G1M+4BeWGcbbSt9ej/wxOZS3z/yKCsfNVEHLFnnQUZ5IzuYukQx
pt0G5nAtUxthr374ARyCMBTm6eZKwpuueyVtzFqgP1IfaSNcO2q42h9/N6Av0FP4KkOA9/iXgjSU
Nfljc5S8ogIGKOgCtz+xSfF6uhfeM2+Z59bf1MK7QVuZyOpiH0WER9CpaNHLvloG4WpdCc3FmcZh
fZJoys/TxIse2hVXu3h1v1RCpI0gqYM44tzGgj0jF9QQM0xqgsjjF6l5QznZKEp09mWR7ZpvOvNx
44poTBJ3ygoqseNDTUAjAjy6b+BNubgC2DDbfFOQTgoC482rGTcI/l9CYukJJtKFOjhpyVyIndqJ
Rw9ZomfNEY3hEopFx6819tnVhfI+/xTqODG2VqSZRz4tCojgqdQNY0YYtNIRb1O4cgl+HXtQ4CiX
WxS3ONEPrPq5WtUkMDGUjQdULonnt1kFekInffPHAy9C5HdGsVnJGbPxYp2QdyWI+Vh93et/X0LX
dGBtjhuUgmYLFoXWG0uY6oubBfgJgD5NUtXkikTJ7vR6G2ZqCX3KsvhCEumO5QZPcpuBzkgrTFe1
gmMCJHV3SudEt0z7KeTgNrK/AclNiKiSUcyWTMRcPY4r8XZGMfsr4NjnBe3ne2c2wcqe3kGTgkNJ
oBpnBAzJLmmaEEecNt4g3WDEZi7pc/A50bU9rVhQFnDl0tmb49Fg0ZpgF8rVJymipggyQH7rtP7q
ZXkHDQFP3ij+dWD8pIkZ1Tw7VKq+Jgh8c9azRq15tJ8zRuCuzDoqaR2PWUWbFLJvh+qCCOP2BOij
jt1hjJt0N++8JpHgoXOgO6/YB2BmZlwS3zVr/AeOwwsUtH3Cmzff7dcsxkmJ9v5ywwXWpgDwPHP/
IVaorzI5Oa41BauURlW0BTWeA83RfZjXIwsHbB2f9Swn3Tou88bs3OZTMxQnkJj0qBh0Q1nngNk9
yqjS7ajNGhVGzsXhWLLfEaD3yzO9VzZ/j1doPkarPt/bwZ8u08Uhct2enC1TIYrMoidTjDRsbfjP
Vz2MDB3Sf2Aftv9zzzvPWs4zi2v37g02kFT6VPqZuib3RNrxCLE+r+0h4YQimsz6MAabmhxvfC1z
RrdC8ckN7thE0djIgTyhYwEVo5PxrjRIVGaT8iXGg9W/eQSkg5tmARkrcyHllHgnirktboA/adj7
LmkHdtzR2n4seFnv6R4ztBFjItGPTtIk9RFDXSmetIv69Nq2p2R6QPZQXNon8y+yFvmACp+PyJnT
xos2uuMvWjCDHnuljDFr5A75it7MNLkIyYEVz4iR0AV9gmVVTG4R04htOxzv0/iDjcfTG566wBQy
VkkzTy1eOppY/k3qJF9HYvrwyE1D57Py4yEUJ42AIpZbkdKj7hO0wUkqUYBTvRhCGyen+vCTPiAk
DwF8jY5haKSWY79AOICFmsfpC43dibGpBPPi1jaCjljh9RyER3t8Brle7/t7t9vqCXJq6EoWTjYc
2j6pGJdaITmFNCjFmDla6tJ+433lCm7u56bmWjHk3/nnrSFtg1oAXFMFg+q8hSLKsfILYUe4Y4ho
2aE6Z6wgp5lKOpV6gylMBisJOhfPkQpIc2DvI8ZI0PKVKcl+ULwXK6zxF7N9e6kwTTRuLYsRmwft
gIt9xHrLPjTsawTI27TObe7XgqI6H9BkkIlVxevXzjuakD9r2QNe19N/3gARCtAMZfUNV7hxP/Pz
FF5PT8roaa9w0dRALHaFBVBAJvQeptiZefT1sbc5la7lzOGkBS4p8t7lZwYiTR1Rsh5/P/HW6tSC
6aeZv/dpCZqIIulbIzYKXZuq21pgzOs2/Mxe8zguPEc04c2FC4FYVVahVNw9Ef4g7kE9Cg8yTQVl
ahQaw549e84no4ay+XoJ2h+AxdAXq0FSpVkPZIAl0udWWKA+JKve4sxeXUb6orUMgtCmvz4LpEOQ
cnYjYVkjeMbch4unfckob5s9JWOdC+B35tc8om5j1NRcND3Cb5ZcaG06a0wh4ViD9ecgowpLc4gf
347AROtVI3zXPCbSV4ad0rJMkulzBIuXquJ5SGGsM8SaxL48zr7bu5X9Vnwf6Am5IUsBOuy2fjs4
z3tmHEBnnmRTHS3jeKh1beOGrS+gCAx9RwaLiUUseHx0imSI0P1OGhNMLA68oiBk1sM6JwCxZEp9
Bzp5mL3Ltuj8dCqhy/FYOQQRRUNjxREBICu2x2Vzp2wlWpg9CO5CSk5z6jOVQB8A1hDNNtQsjeCD
hxPnh0Z+TMPquT7Sxs8sZRwoBKji0SsB7c1XQk65QChiqyVfVUH5pfv90g/jhxSEFN5HQXsBLPi0
AxPuUUAWffQ4iljpk3+R7GXt87BVxjcBlrXHNo/mNK0sUxYV05aQLY70S2DtVmC0o6IsDPmArZcw
4PcnFy2OuYevO4Kl+l10MyEb2RRHvOlkc17agVo+90qL10QRh6t2T4grftIIcaVHmFx4GHWOcIOc
pN1Fgq0buxpdU9Fn/fJ4uh380B98wJZE3TF5NJx63QNPM4vwYFsiiy98bQgkHiM1FT9TrZHHqfBC
0oFXqqubCzxeNE35QZglQ1wXG+ZK5dVdhrYBk1Ywl6FXZ96iJbg9s02BskkrB/i3k1nUHsTfViu8
q7Fi4x8ib2z4CofFZgRZd64dDPlVnOc79IujtuZPnPLURLL/niwMfx5DchniD2qdldvKmxDYCVdZ
dI9xqPndddcMdYmIoOSinJ/i1N+IKjyCRacyFpRB5Gi0vCvvnrFVwrTBwMG/bOL/CI4tvikqWpW/
Mfzeh92V7HnkXJRc2Qx4c4YRRi+ByFcHhiBV9b/fhU/HqECNouE0Wo6SG14Kv8wFsDS7ByKQmXau
351rV8RS9QzRqtut5UuP1iBaE+f1gPklrbbAYwz4AHi/Kc1SMV1KWvxnNkMo6ttLWRUH7sRDC3zr
I/X0LVQmSntWEjoSn7dAQGrjZZA6ins2LWa9tdK7C52kV8cWU1yckEyxNgZjp5Nb5KA2G86YS80d
KnSJM1x2irfVGCSiuxZqlQU/ZphAwnxgXmFoak913N1KRMEfzNTNYmuYQRvOZytreWaGdblF9v6b
xl0/uY/ythPf55XjRVUfE321yuwvHgxgLc74A2zUoOEpSDPzoQERXDWOhWp3E2skcbKfFWtWJPYN
6cWwVQRLNO+3pDN6TNL1l9iH+64acdNL4khCgEditQu0h4/TYhixlAzCLgIqGsF8Ym3LSEbZTbbJ
pCaV4fzJgxCZi4VoERC+8+RowNURA3VOATE2Rjf52lvVz7G/tPH/6dKgAHMV4umvk+gXE74awyDp
pVmmyt5/1m8mEubPGLhNdhr+wNBbzOrpRq0a5uvKJwvWO6i2gfSxT07e+eLrZc3d+zKpHtWSQmrf
9wRHHKK0Z8YHb86Bf/2XTEK6skecRmnO7mn+Iu/MuR1nskD9gmNIYskEMBm9l/SnyTNeGxUYkO7m
tuZua75CqBvDnQTH30qEIgrn62ByQYvxvzSRFsUKEDX5bbPujVdmgrdye2DJpN03Qbpvtb28cKud
XzGHAaE=
`protect end_protected
