��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊SR�5y��R(�*~Ȭ���i��&�@��8��b�֫��e�ܥ�5
����A6���	�ႃ�ZqςN �J�xt��U�ڏ����1�θ%M��a؊�{ #�R#s.^�ҵ�$�6EcQ��:6k�ѭ-#�~j������K��E�%1u����\8�o�UM��攴���~���<ڝ�h)��H[��#�R�����8�
o%�����\�?a���Р���*F�h��b��������0�����F(�����5te'9��0nm���9��ݼ�;���zs�9�)*��.N��W�a�^�\���>����_�0`��^�r4�K^����p7�ݓ��q�N
�ɳ��94�a��{�yꌊ_�m>ѢX���S��a�4�r����e2nilV����k������^�w�y�����n!_z�Y�+�מo9]R@�`��	z*Pr��5S	F7��a�\ރ��j�� ��TX����gnoU�"p��꽠 fmU��Ŭ��N�F�	�u�׻��j���C-���ꇌ�ä�ó�@�6�Ɗ��64�+x�&?Cr�#�>,�:q��>8�s��վ�D���N�]T�n�����0���� �b�X�o(�u�*\���2ޕ򷣯��7j"�N�Kzs6��E"+���ZL�F����{�܀�dL�͖�n�B�f��^�w���ԍK^S���Q!�{K�J�JX���
��خ M|ֱˆ��CU1���������L��]4��t\-�Y��|�@~�T�5��O]�z�N�������%G��]�t�Nv&M(f*RE��!iئ	q
�l�2ׯ)���A�6���2��e�&�uɢ2/��WW�����P�[��ha:(W�n����ӄ��J�Fށƙ�V1�����E9]u>d
 '>������ʎ#D�PwA�ύ!L7pwtW�U����V9}ft
�$�q\�=�o�C$��!T-�0)*��&2+iQ1�kc����Ƹ���N:/������STX�`?�l��v	�"�my������#���	ɩ�(��52#�䥰,IM�E�Gk����]/�NvL�I�4����MإY
�C6�<H�.�51KPBB�YD張T�Pʹ���0 )	�JdN`Fdz����>Ǥ��"Ό�Q��m	��-#�5� ��������yv%g��AD����d��x
�X~.;L'�Ig8z�؟��h�{����1��)�_V��C����J�]�p4�%ݧ�IKP��=\��מz~]��"�F�[������Ũ�,H�Y���7f�V��C��$��;�u;}�]@�K0�����D�����+^׉�����9]�~ȡ����6P�?w3�Cm�*�%Hf��d�)���;�[�B\���B��	P��0�ٛ��W��Ԣ_Ԓ|`<��C^�¨�"�m7Q8����m{c��v�_ʚ14�aM�T�Ձ	^�F���|�5���сE���=GW��I ��~,c�Y�'���2�|n8�Y�xb�_�ި\J�
͌��f���.ϑuo�,h%:s�6��Т3�u���Ag����h��m���>O�u�"fk0$�]w��k���x�ff|�{S��d �q8�L[.Q$Z�3�v0.L-)i��(^Y&雙Q�il�흋d���#1{�T�Q�RK7�c8��9���|��H`�VU���V�LX�8�A)�8o���VZ�?�gH�f�ێ��&�S��G����gN#��&	�F�,�wJˮD�v�>u��woF�溅��[�p�J����$��l���&<�����%�b>���W7|%��7�ꇆ�o�{�F���i�} O���H=C|X��|֩!k��[q��CΚU_���Q�sB2Gc^�B{F�H�|j�Od���Ӓ���v������ ��'H|5Vn��� $�y�[�"e�!`r6��t�OUx���wM$�Sx�,��&]'�]{�F ��~��N�7���R+���,�ؼR���͠��{�O�r^*U旵;(A_$D��������pa����L��38�����*ܾ�fL���L1�v�:�c NϦ�{Y��+Ck=ycɩ�[ir�a<�H�ׁ�=�