-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o7TihX14csMYnunlU2r/PgdmZAnffTQwAgxHz39MucilFvyVkJA7Z7AH5mxPK2NuHaKhk4Ll7azm
NZ+Mf71oTACnKZeCbgqXWrfRNu8wkj6CsjlgIw6s6LwWmGw/r2bJXG7DX2KEZNSsfB/kcXR6y1Rr
oCmrljCEjhpVFIBoMNEJYvlaGtDCeTwG8tFWR9OJn/c4eJLf1QcAw/jpxTCdE3FkYqrlUse7kO94
DV9gxARY5QKVjJg8ERlOIDyOk052KaoLh7utCzL7UmRdqajktkj2tjnb7hoboDoFN6NHzyjF8Gmq
jgGz7sqoJj9HwyS4q2XXGsKorBEF/M4KEYpEFw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7008)
`protect data_block
dKU3V1qPNdsRZ1NH6NY/qJiTuqPD5bjwd4AlPYszNt4L0EfQ+NRWMUxrcq0mVkAxFTAuA4y28+OY
WBDqDdEPiGjjGN74gLI5YVxBFaK00X7GdbmEDT+OGYoJQOHm489CcSn9Z0kbR3VuaMCP54pVTfPJ
xMZY/awWK33OLFGk1yBUYzKTgGUI9E1gNa6LGhtcSCUyxGU7d8p5likczJH2rbzDmKb67bevb7Fa
aDhc3235IsSYjNRyFqVCx9XFzh1fzsrhu80kgoQaZdL0Pssy+twN2wHT8u6YbXXY83aOKVVYDl1W
BrATYEAgEeL9wO+qTMeHEIYFagARN5JWglA68bRmMvl/Xah5BN+Jous/fqxoEoKz4r2WU/AdlAw7
3YpunvM2hpTybrTzoe5UEtW9g4Lx6V0PhQKGNd6pacKO7KwhY7aMirM4Bkv0Z0r/W7XpSO/2b8FS
m/bNYc5jX0/FPV8fNKJGO+40ZTZIdRg+oYAUlVgVBKb0xM4jVlo5twwCSkSoEGRioOs1KqY9Nnoa
YDdP1GBV01V8RRSO906srScS3flksYBzWnSq72bSdVV179feSM0dIMlVFJYBaP1G9JrcfaUrybqz
DGr56l80uIf6JITRHnde5X0RtFYwUyTnJX5VlVLByweWttX8rGsggd7VfjvPDv9PsIs2bb8c4F6A
xHKnwiPe2qKrzka+YPJbro4mP9UddPAoEv405jc0DyIp8PVZGttkl8McSYdnPFuuTI3u76WOziW6
Lec1nSS0tuY1erI/TcAqyhuE7bxoKfYDezcMe9rXPfJGQ1DjdNSptO/TC0lgGq0T7qzEKX+mkWw+
NqFDktwYy3yX5UXMoV56tFnbEiieBZrau9/IEE7nJObZmNVKqjbldATxW9tEzh05olpZ2h5a4Yip
fK0vfxs835yBVLHiKHU8QiA8dnUPc0wgldQK8J+1V/Ym/ZO2H8v+QHVTC6rrfhiTIr3QIH7PIOqL
0VCxNeC/sB7K+aP6MtAWgebR4GPPmGwUXyI/+x+DLSB6b8eYJTGbdkewPZ4VT/hTlX+/L/Db1l3Z
ZGfOsN5UJlOVIC/nKvGLgQR6rNrnpFmGVZyQdPTlz7NII0OfJnN8y6TRXIc9yUKLMZ+nwzK+GxGu
K05Na8hyCFJSc0UygF5inrBqPbwo5bFMC/EkyUkk0SPyU8Wy/X0yncJYnEDgc+GhRDZ5hHpfLycU
qVWaJFXpEtLCIkJGs/mZNdPET4dye38Zf5Atv1cPJoxI3W1yh4uUs0S1rydVF08E8amxQi4KDRIG
DaYuF3cl8V/0oY5z/WOEw8Tx/JGSe5LQqMWhI65j/qYIR76YviW3AQUY/lC0wNxb99HBkgXuA7D6
aafYBzG8VoqjKGx0Ht5ApnJlIjk08Hp8kNldc7cNHNSMpqmK+mlxANi/Ynbm8jbwO5cM2uegpPKI
PuV9IqBqzsuHfiPx7l3RudNwEEJa46+97N+ZD5VI0WEo6E739AVGdq8fPV9sC38IwTNmfAaO+fis
n6YwIB3gVB8ZcXV5PucHXWnBGN571Dy5l1tpYEElgg55RRJvMqdgakG6qRRh4fmx+6pmFFUugCIc
V/kPDrp9HSoRLPSH8U2ilZ8Z9TZKR4vNt5TJE6PSDxeybs6WhbDsjSxd3N1PSnx3BLpEqdjmzDAz
9VvXbTVUpr0o6gO0/4O5A02yiphjBJyh1XpRMMEtWpYSMzmWMhYSuFfl3TL9PolVUh26V+Aa9L//
zViywoJitPxG4Cuaw4FSX8i4l/a7qpw4m6JO8YB9sTWTKUFCVHPhMGIeIRETgxAv2SLEQMBWYAvv
h497s7Rvi4oH5px0tWG1UYjD9IOAMuLut3R2QFuH5+E86y/ArSVU9UMPV4z8JTu2sW1hCaSgVqaY
tl+SMd2L0iQ5mvVyYg3b0pUTN/DXo8SFA4SreU5eP9zZ39fsHQPK6fcaOuUXv4tdAgBicmicWWC2
lqwCCb9idoS+b9FC6Syhqd3AMKY5XU1eIpHyVN3llaFuUi4+4m1s8927yT6rpHJBX9FnuiKVjKVW
96vFk/W6alFmQ8PMQ0aZdRRHYNLgX7bUwqdqhJ3bII3Jna2Q1EADDNvUlhR09SSGeNmhQlKQymXP
ANDIL4uFHddtLmCWeYGAERjZM4pOEqpzzWY8Y/9YxcfW4wPPFe11l5SY8YDv8xeHr42pqZNnFddD
YnRC9xyC/lMicd1LfB4Fsgz/RIPawUW6x9Xb1RTLG9IAEaNedPQd3ezln8scVLBpvZwqvoUFhgCt
R8f52otZVTe1pTC49J53xRF6qAyeqzAMfNSAKKjTWWWNeqxSsZ9wvqfC7gnTXPUQNE6R1ZbHzKYI
bm96c7XQhzHa2pHe1k/UetOZxhFZa3SO7p8ggDn8MunT2tJ8Q4fTxEdHJ2rNB4TGh2IBLtADklsE
6AmE3VaybTnsVbokpq9d+kh4oAx1nrWhPN/912syTfIuTPQwca8zaBu5vvReeiGbb0ymNl7oQ28l
z9YNJykC9yRyMEPTEGY37U23LgN8BVzfb/wk+BEV/ZB4g+DlzHVvOMy/I72X4rU9eB6/O8Z5vV40
OGrFexZ7Pk+mQSLH68eeO6G52xLi9WgQqpHF+V2hxbNOO3k0vpNXQh8cffvIFhWUeNTTkVVikpju
BuvsVFub5qGANQg4rKV1eISsauP+NnTx6I+4Mip762JkCl3v4an1xYeLX/WC+DaFLLNm63LzP5sS
w5fhbOfsyI8nASsCO1WWw+aY3248kIXigS5nyXF5knqEB22eh/XjQHe5gTJ8ks07as6J9Fwvdqas
aswjpBt/wjHfMN63r2Yje5n9tVaW5/Fv+H47AvZ+nsnJYv6GgV8btV/lbE2Q+oCwSmPQ34bjJCBp
NtIpGQkcvOVsQwbjei+XhWX9UNbSvGke2Fmgu7qKtMH/D1oZaQEhnpwSWzBd8TVX1ChEafAixLyZ
Oq2cO0uyZspEM7vldxBS7UpoQcJcf7C9pCnJ+F28Ui8qzjdj6w9VABcXkRUI7qWav7fCkpHO++vw
LSZDNJAfsCf3oGsxxqFqG+rvXTx0N0j39xQf5k/tkWrpgkd8/0gBdSDY/ft3SB96gLkWjxpgByg6
tRx83XhH1SXqAj6l1wDHPaypmR1EeUZQBVcOPLZ++N0Oog5AemALVhuxBf8TJs3WfR2yrlkB+vYC
fku2VLD6ksnJF+AvSsOErLP9LN+0GQlQvuQnWBpWgaht1VMsZJ3rzt+Djw0WFIzyA3DIDbjsv8op
h4t+9yUWTaa1Z8qNSpI7nMHgKV2F5MAfjX8MkW53ot+yiHOm1/uzsoCC7EbIbUqd5nAEYGl5l0r4
dhf6GDNn/fEJe/JOFgBQmmkUBxRgrzjmuz5XVTDPn9I8RJ7SIUQ9iREoBEFVc+JeXctF+XD3sBys
9YH8UiyzHekaNlRBRmGmDpnxv/Vm92hdwKYttTQHUGas1QhL8eUAxJgt49LTOFY4U4iHLq7HDGfb
jNxyoWwQw3RaSSfq6iicO2SdQwKcMyAcWzC6ErI3l0KD2VZyfErvsQg544l715KefnoWD1GEg+cv
scwr5XtkTSeTE64/5/e3ne4qO2eC+oFbPFpZfj5HFTjfojVJYWZJVp57m8DClA/0/VNwr+vkIM8c
df/Bb+lkG8lZbU8fwQMNl4CQ7cKA/k3+NtRUqEEuY1oPHP47C+b6Zn3PlfPZJwq21P51lKJ9YW2D
loJJ0toAc35zbMGw4E+JXspNkhbminSGZWPtiV7jG767JwIVlgfXTV/bbswmnFj6H2tGaxKQusZV
fHqurMShgytw30nQEH7SLUJf8t3FWH1dUc86jCEKCU3xMD6cQBPUcbgmUlG7aRoA2uM9LV2TwKqt
DxWAAk93ZrmagY7q9wbG0fa4UxDWDrE6nDi5sAPNRuKq/lbNQZ2LJ1r7Eeh+RrXNVucvSkSNxJPu
zmCotSnBYJoBbxjtefMqI81JykUFyr782xVUieRqgHkcby2bkx49ekqvt3zOyiL3YP5Dz9dEQFTL
B2D272YRWC9VnzqkPeSXiJ0kVZRz25it6n5xqUU9y02C39jCZENcrcXo2Xk/d3be1Wb7BlKTXEER
+n84ip9isWX9/JKHnX+yVfKUeGVT390f1s0T0FYoOSQuRulUaHfDXRq53kJ9UKaE30MW0IlBiDRI
PJNJS1+piDFLLgmSzbaVcJtmjHoDdnNSaXRE3ZfTGxq2VQM7vwj9Bp5ERegp3ZypvESRhLwlHCpw
vnKEyfeQ7Ywt+DFTnjgFx6nKeG28d09zGNIbbGgTPvPLV/AV/YwN9rbTX8IuwYSrfQOFIdx8hB1A
YUqhlUPdxCE2j+UOtzeiIOMcrYgciNU5TfOkSNCa7TqYWRnfrPkuxQGcY3PfN9RYJHI5cDuqb8pA
oUZzxx/+1LlEUraRCi4HoCYFuiMFmmWpL/bk5CzRJ/Lr64+b8KhsqEurO01XPfeRpXLb5ozcTKUR
eID5+rV+3XYtlyYfk39fFp+64aswDrvfzleyIVVotoF1z/ctdTTqnSi/X+hyqfddrZ60xN0KeXjw
EkhXhlpl8sM8qe6JX1MXZFacTP7GJBySa1SipmkaRV81zpKVkd++aD6CHDJhsf15UD1qXbC302IA
Or8BFV09OpTD4rWCtqozingkVowjnK4OSdgTajqVK/FmvNv+owQlPelHoUf3typiq9/wyZ7MnOEC
Ve4C2wlclZKJohgeJw40T740GXAG+WsORyyh9crGWpuoSom8DfRpeD2820ob9JdeQzAVfkzxhHmA
q3wvuFyp+hfhwojbgqK1tBJdVVwR3UfkL6M+OKjooXl9aeUEsMEYk8N+rmSTIIF4hKsyNUDACINV
FmUBS65A9GkFFIM0aoPQWP4KdUCTGHrQxbHgU/9CaRrw9SRrVGQleUwFeNj5H2vNRWNoSFePXE8a
FUSb2lcfFoPBpeUEKQGvH2Xy0/W0DDKyTa/LP2r8FTUC/irbwNJkViiRBkKIFSC0kFvUwlfyWZ2t
PZgmj4+XZKI8GMOJLC1u4/PcCjnSmfmUpzKZ/hGa7d4ghR98BBPbRazCtIUNDiQyrRJ6LQXoeO1i
3cQ2yMj5Jff3qZtfEd6PSUJAlO3QySfywVP9B5ZBmE6NTox/fJCBs54qqMLgt+SiNx79pdkHgX9v
mhHpoXXFdRBC+DPN/D4Ozz04vo/btEhUZcu7gQL4jcz3FNRg+vBmPfuXIgVvBWMvEqfbakxQk7Lg
swYtkAfqyt0KU0aZF/yQzeE292jwDtk0AOit+ezEdah8jd5ufqRzdmJww2aUpytrH18WAPLve67O
ksL+1La1ue4/OOrV83esNH7DtlExDjejFyBvtGwFpsIXCgdkSJ/tnknPMprfub/USr21PQreFNzR
/2rGq2AKb2yqfuqUCG2e9s3b8xqg3yRkoj8bwKnsLXe2hltmpuwhCAOJIy37LixSZ72/WFUYncqL
wIn2A+lJGzXteWVN5otziX9dKz7aRFlcuUVEwXv/40Ngih/SrcdEnuFhFb8EpzQbKuD5zjjb7Q0T
B6PpZeDOt0WGhfdPcpZYxXTG2O4ddcdQiquWbsFgWtR57HXHMYRwCf7MWjvpMslOQl/986TFAb2l
nJyhxIdG5Q5z62wsmijFXsbCUbEYHANmwrR1hVfdP8JEnvjAtHfm4vX0kf1+QJganadLKtaGARRo
Cp7HEr5EGvwA3psmILAFVmo1U6yG7MV8LNHXvxSBEmKQ1nftY7VKkal4rcXw76Wuuc8IXTAogU69
w/9aD4FHf+k5GwNPCp59ORfYqIXr+iMcfKQGvv4tRU6YYh1zMDIPzrajAlrXBNShxAglTIY/69No
cYUmRodIPOIM1IYjL0XaoBM5VaPBjdn6vNlRZtwqtZJIiO9QiBcoL2LkSxqBxvGtMEZZjiLD4MG7
+OnfaIWgM0o8gOC9CriYZKlBVwXG+l1xTqFPTCRzrPH7CT1GYAqby9n20TDy7VERMrprHTGqTtEL
dyg+fMA0TcMS8kVYUArtck7TplNn6BAhC32N5ctOrlg1+M8/d2LVn05lftzO3pyKl/Q471CVkphP
j+Je9LhNxWk4Dr1b4kqdgL3F13xxLXcwG8mjZqAzaDSiqD0L134JaQe5ykNnsu7W7JlIM/ieDvRa
ZhF7HFOXn57ybnLlvgpGuZXes4AnBq0huTk3dEwjXisx9ge3aUTlI/noqhGQtybrz/loxv0Ykze2
/k4JNFv3NaVY8XCsoyi2xkdZkj/KmthNnirAZgC27ady3N0EZQTs8APXzwH1eHRg4uFufFDcaGUJ
O2h/7LAz3XoXHw+6WI8PXEPXwN6fuYqWv9vF8HR3rxY5/xSe2v0jUIv3MAgrpJNDQW2IT5qFbu7w
ciiskcQWENjo7ptkdtu1T5Ej4iGGRV7abt3ZcJnuMiuFe4TPn2wh7ZVHs8ctJot/v7Z0lcONHgwM
DOBb9jQ7RSeg3QYaUIwQAAnt2s7bbn3/n4WJrnucJjTIj6DHoKFmCvOsCG+HMqoMMcZB2rmxoLlX
oEyYqQAynIqIxrtSnDv3wqnwnOY2hAdcu9GeH3kpD1tA+38RwOnS2VX6CK7r6u5eGPb9J2ENtvqb
gvCrjn6WrKTtv4IssB3uMpSxl8aulgWtxAZPU9vctLj5NhHxB3BBxOCLNoi2Uw4U6jPqW4BSaX0C
bSyt6bNODL914uTS9H8kW7v+DQ43dwwWSaMEQmGCIjPm69pE+v6tqW4fjmiVtn89vKGeuLRpcCvc
IllGqFjoBO0/Z9GG/BuGYLOdo5Z8mbaOUHo8tb9LeJZMmf4FBgCQyrKadVYTjUcp8U7w9DCskgIA
33UnpzEdLl0Dd0unfQeiMyC4bq4n9I+piD54zOmcPt/MdQb0Wwdtx9siyRQ6LY2kyuYglAAiJWSd
YefQyqgjbg/F3Ai8Nj0OiLu9irPEz8NkgYAMQXr1JyMnGE8zuKFddtT3whOj43+eQlBsgD8AEGkt
BuTGNwlRojpi7CDImfParGV7iOZSzVcaKh5mBGoe9BBlfrsK50JLoVT4sSBfODLVLW8F6NVPJpfy
vkVblftuD54jts3uS/ASINgqJM66/effbZ18sLAHuyrVkXlItGTlu50QhZt/4Z7SJr695mZp2AaR
RcOC5VyfHyCT/BUIVSzmVyrYW6RA3Z6OPuvnRjmx+TIa1M8yE09zLUzGQN7XRNexmM2Eh4tCgTnG
XTYZ9ErPj3bbkWZ2UtXZjkawBRlUbTfZ2L731yJMYpFCQFDqIXgpy1rN/2tvcKOoMeqI92fOq43d
IgNRMB8QHiMxrdZevzLzzlPgY8zG8PZaPztN8n34jmFaNdFl10+TwYh7m7PaygBON2QEGXR6djkv
1tC+M0qh408gaBMPPwQszRIF9Xi/Aav3AbrRJt8o9NHpF/BV9Q1lp4hJSW4tT7B9S85j/ywDxJ8c
ta87W46Tqzy8tCTuCLaHBCSQpEPrpxLijXiB8GALD2by+BMM9OB3zqqCpZai9n+eJdSns6RPImu4
/iEca67owZfi/RjkyXbn6GCLIapcJZUglT+IpxPL8OxHrRXCInNgpj69UnQGHC5g2+lDgMYsVLHA
ZxLEvuHYsC7b1b05pKaNdpNAA5o1Jx5juRMOwdTUvAr934De9g7kk+6IZhfekL4c2sWEwgylusuD
haXX1itpxSY9sezN0Qc0zmQis9pI1Xo0WinwcK9BLslYj6eKPowXndb1SF03KYIlQ7+cssuNvtqv
CyBqCgEVZysk/gCFU5RN5dfoLWhFf9M3Lsod/zbyTWcN9t97muMEPad+HPHzOJRgtnXyeAtBJNAU
i7TooY8QaNlp/bdrcLPcLLHzSSmH60OPMd3C4JXL7IfybQnT3jDF/5igwoYhwbCbE5pTbdtYM1Xp
7/Jv0pW/ZtQKj84RDSjeeaJnIGENO+ydpb1HhmrMs6Xb4Tk5HPt6oyzhvw42RCMAedmIGhotb1ff
uiLcPyq9KS/tf5ycvghw7ap9oqbI1Hdt86yn/hkAqfW2yHWguvDkfz+t8TNAHmI1F5grM3fAotep
wGdxfqlyoih8tImigHh1bOhtfVp1W0ZttgG49X9D8NEiUqVXvKzFAGAkzsJMLte1ZNKbpWGWmvAr
hHhgad8wciENSF1eyLIMXRAZUNes3y1dyc/TAGZGakVfcT6D3jVa0gfnAw1rGJzyV8ij964Ov+Ny
Ye+4pVNEueuD455uZUqHapWa8OQsxwyLqwtHQs2Vu3Qwf2cG+mRjDxomDETtSzfUCibZs27WNTWs
2sBqLUdz0k61xLZLuf1mFwsYKyRzmbIHeLJvtrIa+/TFu1gOvLmU9gdul5Okr6s2gdL+4AidZ6g1
bWDLF+HYXEwxNhxRDQZBZJEVXLu09MZM0jmWgeozGLVQNT3h0KGaXu9FWzwZQBGaZmqKIEJNzL2o
CeqTIdkrIzbtDIOPddTzOs1+ATdmrzGZT4nFPZfNdW2M2q6FQyvOIsW5xEQ7xW+zBNyMOraE0W5k
mVymz4pCh8HxmS40k7uh42Y3S/VQalx2/txBV8kxFCZEPAiCuS/Rw3zMogmvgoudbMtAyIuZRzxc
HZSho3b1uGg2NcTVHR9b3cf4433Wek7c12Jn+CaQTXvzM3M916wYofK3aolJniJQaqtg/Grc/55F
GvS1r/2k29WCqP44/amEnytOlCW++1ordvqHyzGIRFtcyCH/0lnwlQWUHKq3AXlrdpl47Q4q3yXR
BUeGl7ONnsvt6RjsKI4itLgmQXbs0NK8haAqRGu+DBUB1XNWK1c18LUrtMqQtYyNdP0a8CcLGrbR
znvxWHc7MthD8ZAUtdj3kBl4qoqakrrUCg8Igmn6lzrc+qx95H8qqY/30t4cSkSiLS7tSrlES7uN
CicFBIAKs8UD0341UDBWVXgmEezo13uQN+YX1ILgu2sLv8L5XKmFnNiiARwj7RR4fd/IGCAm3adq
LcKZ7RC5hvc/6NQrXbbcOWP6uyU9cbC5QTOb8eV/LpGtYhowAMGeZVe930T4+K/7JDuqaszoZb9i
CMuDzRVR1sTo0Hl7KojkKi50JjVGaDJBZWlL7cqytA6zvWkeoqAlYXBmaJ/7NSO5MASwEnDtWbjo
TR1ocbjXg0MINK7ohaZkUlrAdKweU8t1DnJbDLmClXZsHUMswpHywTo8n9V19OFU6MNYfMLfR+Xe
xALiHhOcZpqqbI2fh1fqK5+9VYmeJJqwAJA7Rr1yEQDDPGp3DZk1C9etOuULiWv2ENoy06WK5ozx
Q/qQEhSwn3YRyUlMRubLJGKia2zECu1y8UlYMw9lsEB0e8EToC8FHIxwfqadqpGqkao1oZHg
`protect end_protected
