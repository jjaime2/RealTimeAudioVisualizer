��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���B���Э [$�V|�|��?d[Ѭ�(��7 ;�gG�����h�y(�I��Y\)VYy����Twr�#���e:o;�K7s���b`.���ݙ�%[S&eb�pJ�J/a�Z��W���M�s��&��Γ`:��57��9w}l��Hcؔ�T���M�z�\B���qXb}-�m�E2��W?�.r�0"==�v�%� J���%}@Q�\������Q!��:(�P>��c]�22-}Ъ�������6�m�Ґ`����vb	���׿c0E;{yL�]^�S	�3X�H��=�<�C+��C�M�K���OP���!��\�APŜ}��G�cu��6g��VK�T[�㵒rG?�Ң��:\8kʝ��G���m������,؄vh��;|�4U�mT���*�}���p�d�O,�`�x�oLܨ/zgSw��s�)c;1����=�睍�B� ^'��{��hK'#�1h:�AF��}��m���F�3�����%�%�q�[�J(LoEJYj�H�Zp�\��%p��7U��ˎ'�Zo��j���
�}���ae8T��_����Ht�J�I���Y�Pm��.�O��+1$��ZF'�������A�뱬�Xx��]}���k�������g>�n��K�v{vٞ�ڕ���'��$q��t��bi����E��N���:�i0�Pc���ݲK{�l���=�>���keG���AG�����3dew���������%7�c�'�r��B>��
a����p0��a�fx������te��v����P/7���d�6�"��SK��{	vOM�K�m�d�m,�g�����|�3�	!���Pm�
K1�X�A��1F��}/�*��R��tP;ꄓ2o��)�Ǟ�M���*���jQ����Cu�*��٘�7ӝ�T]a��c�9�B�h�[{P��m�_�J�����
2���D�Ӯ�>u���q����_$��Y�i�}�E뛊��ȠF�\���z4���qtR��Z����^����t|��������О�+o�?������!���U��!j�F5�����#SZFv��ܔR���1ٵ��<r!Ru�R�HͲ�]�	n�� ջL|���P�+w�y�d����|X��N�Kx+��_��j^� �r�4208�*�=�yu|9ֲ_����$�Ʈ�*�BNC�K)E~Ac=������w������`��jΉ��<��r�2^�9wH�z󈊱#s�R�=c�	�Y���1��V3����S{N	q���+hJ����w���r���2���2i��,+��������r�)؊?%�����r� ����Ŝ�~�X���T�!�GC��8A�۠��l]��	��aGN�$�?N�5���~z1�����߂�X�Q;�mt���מ���GT���2V�GQn��w{�[ɗn\L�( HC�І�wf':�y�Gy�K�R��j��9xdY/La�t�Lw��@�W,n��E �{��p�P�
��]��ex..I%�*��g����BP �\<�/�(?��HxC*�Kw�a���F���Q�\��h��J�� ?�p�>'�w��<��SD츦� ie=�*�(F?*t0�ÎgT��(��@�n��'�6鵂�A��p�Y�Eլ��������m8�AV��ص��� $���%]!��-���pFh�Jk������DO̒�y�2��DJTz��[����K:�!��[��N�����.�V����l�{k� \E9�C>��z��2| jH���1Ω�����=Ž!e��1T�f��ʴ]:�`��-S�G�Vd�cְ<Dj��c�I�H":�lm��n~��.a�����b+��^�@��d,]IL�^��j����(�{�tlB����pt	$��좊�����Y�M, ��Pꭳ�H��懑|�����D�mN�ĖP�vy��F��ji��~q�J��x��-\��Ԅn�I��~@�qr�_1�}���z	CR>���Ù�\f|Q!�߾I�	�[]E�0��F����h��am���zj@�lSH�p��J�⹤�H��l_�S�1^BQrcS2f�O����kS�'��T�ʞ��9�*+�T�׎��|��� �f.��n��Kh֣شFݽ;4�g���*��ԥ��m`��؛��,j���64H����VB�D�lcQ���s�j�e������:'$��bc<mE��D쫻�X�Q�+�\���@�Z߶�ؒ�-�<4��9,}��ŕ�k3�v["�2�>���ٰ╉X�b�1�o��E�|:)Mb��	���-�����K�U�����w���Y7j􀤍��1 �@�/}�^B!+��7M+%5��M��,8*�f�U设�L����0@�3�3��l��J�#������ p+��ui*�(�>V�.�x��gb���7�����'@��0�F�v�p.�G�c���5t*(���,i=�pQN�1��]}�Q�2���6<wX�	5��f�q� &��h��� $�%&B2؞uZ��:q�ԞE<0������ ِ��{�mj�wf���;��n�)����d� 7�]2�ì�9������}�k�����Z��&��A'=����{����?U����nN����R�౟�b�;�:��C��p�?\f����n@O=��κV��~��9�JC�
�q!"��}�����Ki&����g�8�z��$�q]%�� �� �g��Uh����&�g1��P��f�L ������`t��F����	O�֬u�9{"��hPg�<Cn�tد׳{��]i�ߍ��%ҥ����'�X���52Y ��|�_�q�%��j~�.��d�C4��������B��t_���-3���ˁ�K�*<8h���!�Eͤ��a+�3#�S��mv��-�&��-]�f9O�#�[�ޟ��d�)���xDQ��|�:;	���I�7�E�]��n�D�3/�4R㴢��N�mӄ��w�HP�ik�8]'�"tW�zx�]�_�T���s�=��h;L�3zmW��Y�]3��FL��R�����<YY�a8��Td��9�20�p�̚�p�ϫ��`��w���0ý~��Ҡ��j�o�Y��NrY�,2M){t����(;Kz5�A��1���{qS�$�%D=�W��ǻ����$x�m4> 1~Qa���ݗR�D� C�Gj�rj}7~h�	w�c�F�Xj��3�����%�Ok7�f~�/�V����䞉�� ͐����v:fR,&�b��,��/���2�3�v�|���g�DT��S|L������P.YR��ӵϾ��^o��\��̻UC���I��a7��K���T�tϧuP�\S��g�K�J���H�J�Uڬ�����FpQ�3���XEh�7���P�q�FֻN���VL��K,;��W.=��T굢�yg�����J�9�����ղ�"�w+f�m�!�M�4�a��P�������ۢ��*�A����D����]���K�����v�f	p��g7Gz���t!����β�BF���'���g'�	�G&��Ȗ��'Ր�.�锪��do��׷��5�&��,ǃ��Jْ��`#X9sV���O?	�� ��?sv���)`�$���pI��:wH~=KS�̾��k���E\����UM�ǅ�l3��kij�mĂ,sn����s>��l�?��f�}��dwAd�磊#�,
�46�:�Bk&�u�qgve��������cF�s�Rݘ���б�-U��K�Ule���]�Ty�|��xJ�/.=wu] + �Mw����A�W�3�צ�㋲^��ܹ�?�%��~N�}7��`��Ss�yV"�d����l6]:�}W�/���ܳ �T��������n��
�cs���Fa,E5�gw⁄�0+��H��s4f�m�s^@9�b'�U�#μ���v:�	��$�k
����(�/���xУ�#PF�it�8ӣb�5��ǯX	/�p�9<���\|([�w����c��[�2_�~���|U^��$L�,�C�3Ij . ����c�ݥ{�/�<&cM���T	-ِ����'�o��0 ��cr�e�r'�A{�mV�\PZ�<2bz�1v��k��8~�3�M�٘.��fY��F��'��"H�Ryj�4e��:s\0���,���4�Ԩֲ��;�C��lU����T���-�:���AFqC������DڙI������;$b
D��ڻ� ��χ7���ƫvÊ��U��=�_Phr&�e���G���>vqbN���ti=������R��D��I1{��J�����C�$ �o)�0��Z��� V�ٮ��=���!�|q���I��4������x�^+q	^~���:��q������5JG�s�X��{�<��#\�&�F�Ӂ|��^:E?(l\9S���p�6�d[J�uG�Hi���;S4�G���}^�
'�����>'��v�T��ӿ���}�F`X��{\�#�j%�nI�xV}�pIS���6j�S��N�c^F�c�d��|-��?��z�w�-Q</NVɁ�"�n2��5���e�5�:<��!A�ʣ���ţ�$���&@��"!K�#&�ËE����)�N�C��?��ҕ�(����ء_��������5`��{w��H ����*ht�Wq���&ud�^8�����|����W��,6]zШγ`e*��8gV	<�&��e�X߉HR���I��/W� /�(���Ǭ��֕��$�q�w�D�&��=�Gf0��n3���ADojB�
c�����b�vV5�����@�lX9��s��=a�vxN׼��n&�+O��@^_r��!F���7��lZ���O= ��X���4@��.�d�Y
��>YlF�d�x���������䃔J4[1I�wøj��M���AE6SaN��@3}쥥$��9������Iӱ�-IO@����� V;�01��?T�y.�^�K.���{����A�Ѿ�j)��b�0DO7�*���A��ݺs�)�o����U�!�����S�� ȷ�sK���(��[݄��w�IL���Ѓ[L�z��L]�_�O��	��/J�,<�T�r�j�ꀮ^�s;��H5&YH~c��m�! �B��?�9�.��R��-O���R�Hz�@-�Lq�1�zyq�&%���
�o���IE��"s��ᇊ�LHh[d�� e7��6?��`�5đ�m��-y
j���>�8�`��f�&!�XD�Q3 � �oS�aF��T;��\� �Y6�Me5>w���"���D��T#�d8���
��`�ch�����Rz,y\���@ѹȖ��B ���<��ˆSm�����J��n6kܯس@7!y,/��؂Q���ʽ�-�39��!�愰���s)�T��g���)���Cᕓ�:/�6+q��ĭbU�ۜ������x�,�ٞ�>�г�;��8�M"�+iP%�x��d�Кn}z�E�!"�<K����A��ۥ
�"�� ���g\Ш2n��D�l��%�@�0R�Q\%I�v\�fh!�s��DA�%���d��k�B���OKk븡�	�$�s��݁��� Y��u�	��_��C�J�����t��r_ܼ{򾋏U���|8{%i4j�*QAm���y����yHz�
�6-qLC�����v0��ϑ���	���EX�kL�Bb�Cl�����څ1�8tI�x�>��o{����-�$c����e1);�.���֎O$��F_j�c.SCw�HC�ׄ�O<�v��Y�T��hz#���m
Q(�6�ʑ���3ɭ�n#(�8J©>��$��	�3�;>|�f��PT^�g53"Q�|�Z��#��:��&�`�I8:���TI@��",����,�����5J5L�R�S]����Ew�AL%ϙ�/�X�`9g��4t�M*��1X��w����^9n����i+]�_8 ?�P Z�/�R �k@�o���V���0�mɃ�!��u�k����;�9��ib.���`��8�+�C��W���*�ݔ%h��L�`@�Γ5bv"FSQ�:HT*��F#�A���Aߛ�Mmy���d@�{�>ަF������$�/��Mm���Z�g"��q!`X���8�s]��������{�U�������stD��z���so�Yq�2�d����.����lg��;w"���9Uu�� 3�/&��]2)�Ȼ$��K�Z3���TJ}�FId5b�6s���W�}cF#0�zaΟ�d��񸪖��@��}'�[�_��gKy.�yT&�c��@"c�'�_|d���.�>f�� �٪��I]aP2i'	*`]��ݼ؄:�ֆ�FY^�x�T��\r��&v�[h�.Vy,���:��3��E�a*a����v<��K�K�HhR�����*���	O��9�'��.;��&	�A���_���~ܴ�x�
D-cb{�X�8�=!@J�3�vK����9NoY�������c� V�u!�A5��> �F/�߈l����/���ݾ���o��d�G\�����
w�_�+���������?W� �k��@�Ϝ�Q�mGW�r�
x����2�W��ȵ�dӡ>P��KһV%������L7�z"��I�GԾ��A���gd�����>��,�:�Z��1i��`�2F�g����%��DaI��g�}Em��	��^�AO����*t��@m�<��9[�-щ<#�9x��*+HqpK� �L"�븽m�5���r�ݪ�bE<e�Bz��GӴ�z��Nΰ����P�K?�"j��$^Q����WJ/T��(hrovU����S��&�7O��_�?�:3��{����]�zdA}U<pY��轍�:��ɃNJw���㕷Z�8MX���I��3��4/���t|0��.��u|��ħٍ���*о�����6�O~;�A���rY1�W�uK�r^ʺ3��sH�f�Ŗ�}d`rA���O���l�%��#���*@*���-��n�QHU�.�d�[�c�UI�ŵ�u�D��6�A
h0�\�w�KX'�Um�����R�A�[�k������04b��4��i'C��ň���2a��@��x�oN�l���*�FR$��c[���.w���s�:��D�_M҈��-<ͥ/2j]�'o�w�%�*j����c�~�(�4�-�^W@��T3ٮ��'~s�-�(���0�� e���"S4���E\F7Aj�ћ�B㈋�B�K�x�����k����7mS@����5>b!t[f��~�p�� d�����]��T}/_�g��܇=�01�9�� ���W�J�S,B�S�,����1�������H�N-B��SH׺��/$��C�nC��D/ @G��ݭ�����4�4�=W�wO��y�$�/�Gp.�i]�b�3e��9�J���h�?zl����(�C�$[%�فt��X�p�
��X��fc�,����Ȼ��AE[�����A9J�h���dȎ�z"XX>�V�w�(�M�Q����~�,��i�L�^�dO�դ$٥\���H٢*p_�7q�
ʮ�k�7u�L]��p�ٺ����<&'ˁ���y�>��{sP���v�!�ǎ�ضS��T_��dՒp��R���zo�v�	5�� jym���z4������n]��%�d��M�q!��o>L򇟋2t��{�i����.�������t��U+��� �%����.D3/Q���~/�J:/�Pū����M]hl�z����G
'n_MDv�٠�@v�.<���|��ϑͱ �Q�������� ���T��B��|���� ���T�Ą���!���P��eIc�%�6��cJ�v��/x��p�IK�*���Kao�O�g*̑�y���&z���Q+��>-<hk]"���6N\��� X|���.��r�Oe�;hS�N�ځ��*R�S��l�MI��+_�.G�2�p��Rp��1�&�zy���YB���{���Lj�x�I��rK!bc�X��/���9riG�,��pn娵�Y�lR�ht�
�cE`�eH��,�c+�7�d;�?j�b�fٽE�`�p��x�C��&aP3�V�Lr~�%{\���~~�]���b^r[���?ӷ��]�s�g>�%�h<@2��|���)t@K�>�F�p�t��G�&�9S�t��Z�^.$7W��D_��`nԬl�b+��l���&�ލ���]j 0��A}�>��.a�Z��z��J��&�4�D|���C�.肇�W�.���tt�����1�DVLn�+������U�ӥ����s]9 %l�ρ#��
�����:j��t�������\�c% !:��C�_�b����U^�w@�i��dXUCB{\��	ߊjZ�>0���τZ?�n��0�_�u�s#�/_���Ga�q�Tվʢ�8��ve�����+\��F�eѫ"�!/���,Ң<��M���t2�q���8�͐Ba�T�ͤ���`�c��O�r�[Un� S�g�r'K���{r�����y__�y���j8P>fg{�x)
d����� �He��X4����h��}���Xʦt��X�RL�O
���n7����j�%��C}��\����y�;?��.�Yf2}%Ǖ`QT�پâ9�7�C--t��2��!w��`�~��"j�o�$^7M��t�?"B����ǐ\5�t0�$!s6���K,JJ�Oʋ�݊��p���.��]Oy�6^�k�I���J�N>{��!Ue�8�c!�x�?��,����)Jo �w�I�韐������:S?Խ��Q�\!�`�wX�����Υ{<��w�a��S '*�j�==�'��Qk
;� 7�p�X�L�4O:.Ӯ�0�U�ӳ#1h>��M�L���{+fgɅ{�b�A���2�T5��Ŏ������
Łg���عb��e
:F�@\��~X�Yh�X4.%E5�-x����mJ�\��_��z%�q�>�1�V�2"�rY���t��ӹ'�!Z*�&�g��P"��S�^�0��t٘X�-��
��	��������\�-5����9�@�7dL��馞���F��}��w�T���(�`�o�xE�.��X�B/G6~��%��s��s�ػ�M{����acۦ25���pF��{���齡V,1_\_~��pAA�|�8��/�^O�ɠǜ��X��~��4g�#����Yj�-���f���\6�3mH � �v��1�B`!�('�r��q��0��7����7����@�Q� ���XH��w�T���!U��w����Q���,��K"��^�l��˹���3�+��*����*��Kʺy7װ1=�l[�b��vs?�{��=��m��~�Lg���|�y��fĢO�M{�\R�`aG=�4Gi�$[�ۦ��G�������g�T�"p���~�/�:b�ISB�6l5������{�uK��6�+K,�����!+�P���ȁ*����3�I'�.]��xKM����kҙ��Q���R�	��)����ʾ��b��靥ʱL� F���<Y ��U����<û1�!y��Ϲ� Q���+��H�2#:jA8���_���n���q�O3���k�s�;����+>%��Ag��&8�9*/޷�"0�E�Ep�}zB_�|�D���ߙ{u�^k��_I��.S��7 x�	�2iߛa�V��V¥y�KC��<�
P�~�1mr���Ʉ��O#��Ĝ���GZqw���T�ax6�fsԮ�X6�?�^���TG������}f)�g��!�op�,C��5�vO�Ҹ�S�gvu�5��j�{?��9#���3�iw�wZVP��:�p�Z�%���Pt�2���i`���U��vqpo�K:��X��h:���`'�O�v�Md����]Z��ΡY~ �ܶ�u}�ׄ}���E�'ܭ}'@`��.������lGW���)��DN���0i�I�H�7>3�N�իp�6i��h��co�7.�R�25�� ���>^SݚT�g��d^��x�H�����j���t˓���kt���.;\��N���	�@VaxM��5�x䓞<l�H��r��]m�,Nq�C~�^P�k��m?=ώ���;4�6��U�S��EA�j��8��,QW,N�>�z�6^����29a��L$?뒞�����;�'R]��X�d+g��� �]�&����:������X�$�/���j��qf�[W�)�EB���s8�i�c��~hR�^�5�
�JJ������/h�I���G�w�ado�j�r[��JV�hO1,vթo���'I��s7��V�Q/�����,��R��o�{j�FSn=�L@Ĭzk��͵W�r�0C����J�[%��1{j�a怍��K+K|�x�}�яΟr�Zv�U��U�k=UZ(�a�soYa��I0C0�f�/GS(f���e�Y�I"E%g)�O��<���-�E�gk!�Ky4�΋�,�,x`�C詶�KZ������L\Ľ��sh�C���&C����t�D�8�BlZz�����H��^PK�C'��O��sOsY�K}(��V�dz�O����A�y�z��F�}a]&�]`WK��K��Ff�J��a�˗|�#�蜋#�hQ��\����Fb'w5@� �k���'\�0`�wu���6s���L�($��{f�0�=G�bmۮ���Jl@�	Ȉ�{��'�3�\�����-�d2��ٙ!R�q��Z0���b��^/��-�Gm��b�E�h�]DB���"z�,w���|�rW�#W�+s�c���3x�l1E�yʇBe����j_����e}_��	���Aʥ��������j߾���W�h�&-T�k�@:
��;��)��:�E`e�s�K�b&�
0A��N�J����D�F���q3#w�kg��S��#�	/>�ٞ/?4�!I���]��
I��P�1��IC�:��/��Ὧ����Xj�ja��Bt}d$�.;�nH�#}w"��5
�A��Ej+��A��6cΚ���U8'���8̊��'�&�ċ�t4Ǡ�p��<(i�o�|�z���'t��M(.����B�M�r�:g�&��~胄d��gA��B���c�-�<g�R��6+B�ۏ9�d~��#0�'�x݊��,��0��N�XNᣄ�
C��l̸!?��VzAת�4��Ÿ޺���t�� W�'�1��w���[�Gآ$��~z�ٟv��Ԧ*�rG��J'�]��yLt~�>��dB�J��L��iK��Kc�Ϥhq���^0�
�^��gCB4j���wБ�n8-�����O9�p5*f	�u%�&ګ��|�u>u�&�ܻ��7sd���a��Zx]��)0q��Q9�G)�Zi�VQ̃�ǚ�>l ^�^�U\ܝU��ަ�
��H0Ѳ#X�W�M�?�*�+ �>�}�|>����Y�-��?���ɬ��Z/���X�?U�8"�M�\ӊun_���0v��ڭ��2���mUqV�l��vn��2��MJ��ta���*#Ǿ�wv�ы�3fVZBL^��Ebk}���~ntm� (�v�/�����ԉ�/�8�%��U�ի��f����/��Z]��?�ܚ���+{34;��dѡS�N�][����3�-�Όʖ�Z��q!I�1s5t�6jYM�������Q�)[�2��<�b���8����bp��&-�h��Н9����A0�R����Z9����0�1�~��(1)���֪c2�p�_�ߐ���G����SM֌	dڿK�`��v�c����O�~���l���,]2I�%&k�|/r^����"�0:�@���f8�3��{_�B�#$�F�.X���*�d�X߽
@��i�g���������"r�}�C����Z�4GwfM���O�ÚZ����htO�J�NF5-��l1/��ETɅx-4[�hB+_��[ݕ��n�d9��
�Y�&��}� B���V�NޭXG:�:з���3�8D}~��+\��3$��b��Y�g�W���<|�A��݋�\���І��l��Mi�a��#�\�n�R-��	X��	����	z�[����Zwj�L��(�!艽�2�����>,��a��.�� �Qܱ��J��e��F�
�5�t���\��$��V@)Yyd	�מcģ���:�3���l��2*��oP�jƙJI�}���1z@����ОyIx�0p󞻊r���]�}zr����r;�4�����X�������t�'9>mP�D�!%� y�%�T(�]�.���NbN#anY�m�F�ˇC"�ܩ(�b"�N��n��eG��R0n����&��)Y��*�h��Ǳ}Ɯ�	ʩĂCl2�zd�)C�;��j������E�g��l)Mi�����er��������/�x�s��H�`�Q��?x�ėFwvn#��aG���c�5?` cW"��G	� �R}�uD�$�-`�I��	�