-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ehGwe52+WAWuPCdFdyFN5YGP8H/QpgblpT9wTWQaYhTY03ARWudTx6ASdnL7E7yawqHRhRh+pKeQ
X+j/isUeWIQkHsmhQdATCDpQO0LxF4m5cLiFHrV/Y10qxF2/GBrnsqrKhvDlqOkO4XE2e5D2V201
6gF875bxrXkxcOzjTKYXFilA7H1ELiZjndS32v819wk6ygyvAHm/bfK0N8KrN3QHUqCgyo1Uast1
1AvItMnTg1LHLUNLbWncjPXizWhHq/3JE2XCtB6yEacJfoL7uTVM9f02E9qYnPPLCbDZvm90cI5Q
tC9jqUuTxCyn651qEzX3tSVk6ihplUCuV+ECiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51056)
`protect data_block
kLKzDSKU7MLKfd7vx9TpRTEZ3iOEYCIVIGe+VnpXw73+/2AxcmS3r8RZIppjMSRokQGZidXsaXsD
e+EgouZyZGi/UApIwp6ud7lS0Z3RsSmKFYJdVF1EPyyUHFHVyyaBGmeLAb4ZV7yAC7HFFDWr5rTv
70VL/fZ6+WzowqhvwLNyzGYbLZEbwEWi8M3MnX1r/fmzXC8kcW6KZMH0MuZIVjo60zlom4ZJkbrs
0NmaZOIg/KlXY5UX8SN71uOVZrQWO5uP2SJ6z9Uj3hlFICxMMqmTonxCIwPhJEEq4iZx4MiHNkS3
src/ZeuUkBj4yXF+UMGA1S/x0C+U5rGZNQK/vBFMaU2kETYcjSEywfrzpa+uoToUwTzpYX1baNQ6
HPxIOVSA3MNnIk8rEsp37TZDj9NiDT3mKXFhM6VDkNn+dikI0S0W/3JJoQruDwmCAI59mo9CT8Gq
VAJMqgr3QET4X7t85rULyXc4n0UVpQK/3lwIfyx3CEraw0bZnlJnVvgx2fkVQ3HSZgeoySc3kys/
AN8L87I9Pz9oAeC9utrE0kIlVI3iqkuy4DIMZD6j2jfuKIiNWci9fHSshzbwllgeoj2ARhP5cs/S
LeYZ9AGFMmUxL+TqSBOrCG9Z+8R0c0TQSiFkjNRu+NslQpyD6vsDoLdzMIkiZrCOUhLl08kZaBOc
Lp00A0o9MdlcQzMQOeysahJuZmaIbFVKgHLeSLUL4l91dlvgcMSTzSOSE57asPK7b0WOUk0/s/Lu
ZqgCXzst3WpO+aPfefhTbhDzrpc8lTmYqLQb3SZ5Ro4l+4muObrkO70NaNIb1xTZusUBNvaNXG5u
BRN2/NBikmO/Gbq2sIp45yfQkN+jViGSe6Eom5g2OtcKKySb+2NLZqyFuo7zZ+urM9PRBSouNG1c
sYqn0O0/GK9FoYM+ETDr5DbIPq+4uTDfWuSSzXqnffkzbwyak8gphuvwL0UrmfWeSinAZqyyHGgQ
cTKcDuNN1AcuCShQ5Bbjxv1dVubk673Y6ID+2Kcb2yscZSZTsJOradQGG/IcK//zJwaVQYrnHgBP
JQmGcwXFeM6kBXaz0d/T3CcIKY2vyVs9puGDputlXgXqXtEhwpfLY30rcms4ZRmb6ZwV7lmV+8Ys
/TbxeRwBkFWUHBq7wXgMHJDmECps+Vb01p6QdtSl26quFIy0XPNByLgN20cJJHKmzzBmW4SulYtd
R1WsT1gNjEYYhSyJGeMJvoLoxa5khBgGE/rLBCokH2yO1fzfd5Cnz7U312uC2DL3N83JLxTMQXBL
kclP50Edpta95+/txWys1bByUfvh+jzndTIHo9OlzqP9Z24EohxIk+v8zBG1ZjMYB7DEm3ge4asD
H4oP8v0foIkKDfDWgE+3jqvVZts3vMrJDXUOg4/Bo1PrYecZ4NQzV+msPbppiHbYS5qH2eovXtlq
4kwOJ+ybqj/idRjW0N7PASfWnMVmATg9Nf5BsKZ7pfQLmAFsM6MfOKqzu/KpOQcCwmAtvs9OwJ2u
YJAAf0YevL79ev7IStMVNZmvBuRQiITuYols7dgEZCtKmReNJUn/axEE2KZRfi42PQ13pbEz6R/U
4qYbKas6+M5r3H96F4SGm+xDKjk+If7hAnBh9WDpJD89ZF+TlBoRvJasN/fIm+lNrAeVoYgM/tAP
KGRL6bpJ8OYisIlhLxOV0q4tz0wUpFaZbkhfTeFl9LMu5aP8iUzTQTT9JxzpxNmkPoC7eVV306s8
UxFE/Uk2i4WEiwvjybU6WO9Z4nz5kffh2LJbKYHRFFzklA7z6PaZmcP9x4uuDGnWu9kYoR2bkF73
P0padKZ3P/0cHuMKvc3JSZcmEt/HsJu61pdXR9awbV6q/rnNU0xbNpF2ai+S86dQM9xj+GfRZLSs
hQJ2RJ8DD9wViyrti58MVusU17Wmv+naYUGPqY/zZnJwOazs0MK7fkGEktqnyXi+qlpYQ0+Ap6MA
LXoBkuLx6iI34FhozwAtjeMY9WyGJV4Xu2obbXFphgVvbsmHHmRgk78bpl4AJzzyqlMAycn3Rym0
64wYgSHTdIYrvHPaVmbI/86M396KjxW+7hjhQfuwTLkgtQgIZ1t4DDnlMlmLhGqa4z8350rcGqkn
uiZuzeePV1UEN6qO0Xp6TGO8YnelxD0G4OnJxE3gTXEjigxoDjXlQ3WNBjSCLft/r3OIdgMDYXZK
WZGPXnxskydIQrT1KIvuDYOWOPrKifcE/D+WMYh7hz+06vW6EZP/T/ptFtS5icOCHmq622izNNjI
xHb08ORGxxeDuYEMydO+zTtveo+PwvLSaUDAE9WGsz45pknMLNs+kYtAKu/LmpRmqD5kJFX+NNCQ
G5jhcAN2QByT6HbsYozF8yn6rvmwaoKl1KX6DhDAt9nwlkF/sj4vyGRYjhgkfSLOe3PoMR06wdcy
saE8hu5tPwTr1LrIRU2Id/yFbP4vGCwnKGWEdy0zjEv4FImuwUTzpW588sCZOpINLTICPJZOpRa9
YWoIV5G9Dhx3EZrv+HTJV3FAj6mWl2PPw/spTGh37TpeVo6JgfU63+c4/hCvk+Ls1Xvb8X0u3d0t
MLDtvFQP2qP7PLQS64RyDu9ClKMYSJC+w28HQr2pBdYQfNr+bQ/0drOcjImDDA2ArLwQ7vAM6yce
PCw2muLOZ4+gNtCCSZFXBkj87RYjvKjmNESZBJ5dYNcL84Kket9+YcADep2hf+BGU4rCoD7s2iU5
Wxzxbmvw9mGIrlqmGCi7P3x9HsGBggzdUqyNJAQJ/I3Bsk+em+1f+31Kzv5OKOk9qRroPCBa7CHf
weIdB9utMgjWHqMD7qZ8QQxr09vm4ejEeGpKMTGYL6mhd2uhTJQkXJxFAtyQLmlQsqbrGKbEoQt0
RPfoUNRHNYl3UZ3/FQvQ6b2Pzey1kSlmZ2QuZ4obJObEfyhKizPtwvFx5h6ClHH8frMhYeUfiTqN
s58AMJD4dSMP/m5s5mNDYAMw911C/vqWEuRiP78YGi5MTrdlVhAHzE5N0KZliZx4swMdryHsLnZ4
vvVIM0/ZdfiVFZodNHA2x9k1OAhYUQnLAc7KJ6WsVyagqVdgEqYeXFgMpjrH/7Ixy0emk/DqXJ7V
dVJHUz4ASKaFBqoM0JOg0Mv26zFQ6U7qiLewkH2HxCxKdgYgiCxD/15HfF1yDH7/UUvL++Rui7ED
FNgN72i3uI+WAzJaETc1/r4F70eYmNM3eLYInDEQaEvudPhSXLjftZNUIcs7I16j0fexs0+dguk1
uLrl+Lcht0n0g5+UBPVmAqSI1voDnjXmPbh/w3oVKUaijukRZptnTfP2ytHpt2w8LFd0Cew0QXYp
riY8x47s1XIKa0z1rwV1DasA/mLNbkrcRgWehxg40elYR+aWcW0GSYAE5TVp8986juBmxwTycXa4
Sop0nx0bM1W50StMzN64X08cWxkjPHqhnkjADne7XK8g3Mgd/ilAcVQ7C2h3guQHZ1Ys6BESYnSE
8FHcue6k19X1iverNspfsdoPq18vTx8VjlG10a32a15BRFzPCXb43X4k6gTLYb8ud5Sct2357oRK
Uj1PA2Xm7Rehe7fI5xvOVTMo1uNWZuP6lucHxoZZ8y6c1+xTwiq1GMoP0WLKbtF2otOTeGVkj96C
NRUbPGYDR0QXvrc5YEnwxa7UIpD09seTN6DCXBf13bpjYUIqYcjfZ3IBuhAnlsKEPmiW2pvnXcIm
XtoC5czHa9xDp5t7mhnyMY90Mm+tkOt3B0kPMEzdsl4dYOSEF7aYt9mfDcD5Q6MR1Oywz9ZQM0ae
bEEdtc7LfBxbLpJCi7KPHU4VGwI0N0pMpCc5H4B8PGZcHJTPQT9b3eT4V2/ppRZvWAH1fxh1y17N
JADZpjU8J7MucK2P4FiFl0kl/LfuDxa4U8lWwH2iKwGcmESM6A93wDgUPCAtCy+HOAPYDgYswhRV
bJI3T3qAuOd0Wj4a8bF8DGpXqdGHZZYRk12qX9btJEbvBd5C6tyztEhWy+beWMziOn1wjT6Zlcr+
kTgyspizAWUqPxBqNx13FFjuEkHg9FRvhP43FAklet3H4quCE90OC1z9UMHiqiVWNNjspkjxDqcM
9ssvcIB/+0W9pc21wf56jNy38AjUgrgGCp6BMEVYDblamVwTm5YqlYElUbiaKPEPctjV57lI9X/V
jPD+pvHnOOCsDcsF4TkAvGB6crC4B0Ei0kQ8+5V/CAJhleytAjJv0lUGajyJPCbjih6Rt21LpHZX
7oebGEiVn+tYCKiSCc7BG1GeUsOx2QQSZUqVVGar1yk+JzRmK9Z8HU4FeHwpwoNtNLL+CbvEvGbt
d1QYbfN7gamE+qLmNXKszbD2qtZkfOyOTO3CSE8OmPckhwYCZ3arOjUICdfGmAHSibxaVAkmNXVt
qluxrFFFIhj+vAc8ioWAzdGiml4DKJ3iJ+iOd/6eY5GvCuCkxpW4ylrj6LMTufmL0RIS2dn8gM3G
x7MaxKAPWmdFQXhzUCkBKNCHFLUjItZMuEQzku98/W2g8vzZlKUOepBAvZMPs6b/bBe7KqyCJLZw
a3BcRQsqF085fuWhg2g/svYhtx3BNVVlMbKlS4+JM0I2a+78nHq/BeiTno+EeFNY+fp2RhVvH4S5
gv/L2tZtzX1NIUw1kng7UHU0SNEQDKWuJZi7JU8orV/DUAJ76tYPERWQdm/Z+50CYz3klV7GKq7G
TSuvUSSDM6BxO6O/DqxcxzaN2S+MwDlWnM/pRbqXUpsij8PfOCcfsOJlZlDFS2jejheoZPcdCZjs
EPNjXPYjC9Qy4PvYZCdCwEADR9pJczvtLyZrEubPZeT6f/QFRe8CQYBqrldXxyZjrc67oCi+FjoX
2C6XlwfLnOrpLGXiq8qfbCluSwFk2yEcGGiWrHJfe1ErjPW2vzfKrXtbcIUytVyLrtvhKG1gAUAl
enEBjhpZXsR84wuAgQyREukRO9+iUtzKYJ/icYMQQ0QT3zMAe+H5E+CsoTtQKiY4e5S6AQyegPDF
ZGLsk3Re0BWEYS49JosCa34IwGx0VZwQJIo4ZMiNAawe4ipcOH93fX7EG/vLV2ZyLXZbJwXs8ysb
f5UjQlQr08Gw08VT9W9yld7aTjJITWKoDcLytksi1gRwL5w28eZ1e5CPVHh8mGyYVOlXIP+FMqWt
XMQ2mgJeuDO2pRYky/Q8onozb1UP7FRMsU81jcSThKjB24XmJwIJIgAEs38PcOvnpnOp+RA7bceD
pem2NVvOvSNFh4Fv/PRmIUUYdvEx98/vFWgpev8EOOV1lxs6CSOsE265EBFWecNgW2fpd7Un0rf7
mwbHpjQvM1fhS4uVpwyWD/heIzflE2rHRGeoxGutG5yYqOs6zMA0OgeSIfEEcETR74Okfu+CkTix
vqjeOy1PHDzVI5zD5i/edp+Fvo4ZWyW7v3YjPXa0EvnZ16CeQn3mRcNsXuaKafZ11WPs56C8ZRNB
DPOQNgcQAlTZiyVAoZFvoDdTbmqJjZKnCMnRJg2bRTyccataLboP1y8xWdN8EU3tsT/5gAFNPw60
pEYBgWTFlHACx2oI7ZvwE0Xi2Fel28+A4ogS2NZqUDT33Qwt85zexlogqQraPYeG2jhezJpzyyN4
XC4gLlUvjJ2H2WCwWKbL3PPYWMWulREb3ePQ353b4sqSWjbEbL+NRvZ3jsuq2rnHonuUwov14jV5
fxTkK146jM0e9wf42wRuKSUfVtGZSczMEtZSLbeJZyntGGJHP8mzlFejhmfVE8A2Utx04ZR3vMf2
Tpjk2zPMogmtLtnSysRv0AXUEM7NO13RD5Od5EJufhRdERomUd5Nq97DU/TioaXvo9lIn+/spvWF
KyqMaCpd/bZ+s3DlySM0dJEPFIUkO6tPjtnTElJGWZtdiqUgcwjSLEwdNVCW5L9TEJ+UqGZ1k42d
Npy4rSNQI+LB8qFf+zCsoahG29kLT1zmyFsH75sBG7annjIObO5md7ZZR1vC3rItWgLBN/nexejn
xZcYeyqeVUy9ZuzqUOTlrjzQnHHS2/Uxatosq+mt+AY4wjNMLBSmd6HBfyMkYiQ+VGvxt78BA/Qt
sDUsAftMR4drgzsDs+Q7/EIQuSTnedwsQ77R8+Hy1xbCahO5+DeLve9G1CsP1GT7mHActrqQWAUr
o09xakdYgPZHMlmmoxVpLG3W2Pa2le2oH46c23tobwaA1nuOkxiSA4fWBZ37Kvf21DAW6t4SgUzE
hhmbJg9jcnOqDs3sNpuE/9LtaD2tqwes4RKimXK0OkdwWuoARxqrnA87z/m0wBMXRjQt87W6JqrE
fe7DcU9iqArutksoQWE4ZJ8rid5+Kki8+eTglYVFG4zkAv2YyC4vFaTv8E0o2mF40+6VF9jPsQiV
p45MPWIJl6QjVrSG4ceq9mAD6F0vE+g3i+IK+gkhZm0j6e8+DcbpEMnkMsU0sZMB2sWgmdYrDpjg
zb3KXMJ6F822it3dSUuKXFHb4UMqwbiSMXTksS/i0s0fWpx83w3NsWxi9eFo0x5D8bYH0j6K1e38
KjkycPDLQGhAuyHaAiYYkkEwjHLUOTPBB5w0HUUe4/Tu4bqqwXZ/2PCb6CLbSr0DTxqrGADCAfBV
gGVrBlNmKk2Z7Q0uGh9p1cxnxPZUMdJcTOqhA531h0Cu8/FL57VrAEJsOWe7svzoMYLLt6Q3K8HM
RB+lUN3zlgZ01tDYV9JrIdjsgEERxHjZ047ckXT7pX1vD9ci5MpZdGTb3fj9PdP6shkzIoKh4rOs
Ch7SRUqJqZcHLD9/ZAzJgKu2ai79Nm642u4dhvUlnNKlNTVDn/durhoGwHw28l9vM551BF06e7xi
pO9Pob6A9JPdWloVgKbcvp9liI7gCSgKpoVI3SxF8jZGl/U3iUtT+hy8j7IrzGw/qRiukOQ7sinI
gR/FyMuQlLHMHdtDIMhu4dkVdud2U+ks0jQcOrnG96cRnvPdr4gUFt35g2qWgMxKm5rz57kl/vXT
s/WGkm+PsmeISV089WPuHRIVNzLteIncWEaU0AtuzkLNgGlWm4CUxRkIEau7CYYqujq1bNxYSV5T
JoF9sREn4qghDx2ZAqEoNbF0z+ajA+dPeVm8keOU+ZcQ1EiNt/GjtslngaSJihlS1XKeyXWQarXE
xQLdkS0jBEpXmoYytNa+/uQzYkL3bLEq46B0AG3Awxa/t6QPlmVoUAl8k5SIKoSFKJSQYtayoFEf
mj3AZCir5ROHXVfBc8/wnxWWPaTJVFlp6YFhWYK7rXdaNCzgqphhY381AC1afQAB6TGhRNhNpwAN
st2y63K1niQZp9CiRMYqpCAh30+ejhVxebnh7CW5iWGM8t+vQVmGcFQBajsshD7ssxSCnNE5ZjL7
8iepQnK+3xhYYaWMdHHUmMdoC4ij8wQGQHXuubY0p6ATrOf0ml5jGu3TlKD2JXoGsFgDSY+LNeVI
hsCTUX4GJ0IQpBvyEP+jpRuTjzkE08s88mQABeIiDgx0939ka8xLfcLoOd0PQwy6T23Rv48LZf3t
NF6wa5sk7g4boHp3LluHw9AS4jlW3kl3OTtwIx8aG4tgZ3Jg/lApoTDskc6R+4BvW/+qQKTVHoh2
OvpX9Ws3rwY16XOtHhA6fRJQD/Z7IxlT5HczNS6S6ikrnGwebmcoGRY9QgQGKYcfhsQ64MP4dYfh
m10Bgd0YYv4NE9TQJ8Rj25X+KlE2TmQR0PaYLP6KU4t0udCb07y7fj1G+P+u+h9uwpONdpNo71At
xRqzXYcappPgbFfcyH2/FBME2wsrz6deFHJLdghwlwdLN7tTv8J8JeFqu7vB5+pXzsuNSq0X/7nc
H3WennyjS8JGdC5tUm5jA7gGE1TtLNP+xdjvs6azmR1rm3TGEPGn9HdkPQx5zvomxoaWa7f86RYy
qntStWRN4Zw+K7F6kPlDsSc5tsnhXZO8mpW4if/wrpDQzyoFOhk02l2qsPsVnLTVuHkq9nBRr39Q
sknXSAS4alUiJ3BiOgrhqgzsT6GfIFIa41RnYrKbBSKIjbwty/VgJPbnQxXnuz9FaQO5KeX7ugOx
0/XttTtNPD/8/dY0V8rAosA/8w6DAikD0MbLEvYHhmDiAhyiTV8Hwf2vk3MjmP2h/KGDOfuUheCx
Z+LADqM6+zyC4Le/sqvSdR30+7O0OhUFWTDHMVHRsyCaRd1rlJrE1VPGjlDH4swuJamCnlKCF3r3
ZBSYJwJesGP4vLTG/I6RvNYwJHHXaIHuf3Xv0evPnhp5XEyoq4NBl70DlQv4qrtji4UIYsqC+4ng
Xgnpdc0rboz46VIxBzUvV1i7PEQid64AUPnEJOo4zXw/jze0M3lJ5/0PHMFPAryqgFvrMcmlFKy2
Z2ODp/+IlsdEPt+KrNplMy88BMRJ80pvgG1Pp9l/kPciP89Y2rsz09q4Y4Pjxzm62Lz8X9hJWc7X
PUsGnCtgglOaegXQzdaticmWjjNacMidYPL9sqHas3VytZxulQrrVyot9+Gng8Ph8pKhSAPPAQY1
7IcyO4jBu3Ce89e9ht9DAhovYTvhi7RrldyCKxyLkHTjAIuPdTwuA12ED1KnprH30nAas36tVxBu
zSPwEXk7QPJWT9rrZoTnvSY1FX2VUKhJ1eBVb9pssZSHQrEXwtYOIJjFIUv3TywaZgFhvey1I+Mo
oSS4QHoXRDgCNvNbDFacm9NEKXAMISxCby7vbEaAxd/MvuQQrZv3a4HE4juEu+d4j8/UfX0wOpuz
e9ZSoLElw2jmGmn79QHywecB721XgdbXxVLlLQV15Qlc+JdczTSSRfHEloXXGzAVMKe0XIriu8wT
bGeinAI9Kl7SvYulVphkEgZAMHtHa0pwv/wVFR/8X2wCsYTWLPQ09LsOXkwEeTWpJTKqK8oSvYHS
nf7KTeTbfVo+NDDd/5mQEeMlC6aPTz7lspK/1LHp9yKN+MUO1sC6hbawIl61EjySNSCjowSbctrg
wg6bTG9H7SGRoMO16ktBUzqzf7bp/Oqyb2n49cGNcC2Ip60rZnEzK3BMrNFC70EXs6Yh8fu0N3L1
bg205wRH3uPS7pLazDrTahlXRcscinWq1ttVMBIpfIEMP4ASYUMnAsecjDP4ODAgsoBsJJKC8hFH
XiBO0vZeJj/jSPZBauQIccvN67oaIlCbEtolfvh0RYGzyIReQTV1D3bNjoas9yrrbZZpGwaOy8Mw
/dnCz55ujnCtDq94Bijg2JfAAtEn3Z0/cQIdzQkg2ab/omvb3F1+WOBizKdH4VkocVpa1lHU7MGb
fjAUX0UJ8kAhAkH8kp+sB9Xq5ehYNZuA34oBHaSkZtZ+/9yJHLBvpy0EaAhFjFDlqOD+SqgJQQcB
Jaidb5OvP8CkIPRsXshtkEo7SPE/Jz0nAtD4wjrIuuFD0NTTtSsrrgEgedtREJWyCmj2ETlJJGS8
7tFYEnFhlOoefZfWO7SeF7y3ELP2bIYHpOAB9h/q5GKl5clsoJSaWshXYChy9cqPCSQCTNSAaQJr
PZMAqF0HhfPUq/K+vxH6O19wzFMrbcMtr/H9waFQ3adExlG3lU4fQ3IKEsMKI57jEsIb69SN8hVU
3xF6eWwzdpm4G0mfJdRUb8Oc9FEZqB8OJSAgnUUDIpHLtbUAJIy3HAh+dOka+Q8RYBp5C/VxPHj0
qNGtpjwsCzDBCNll6sQW3YwaYf+m5mVFM5nC27Ny8UZ30keWV6aoXJEB7wXv5BqGm/rh308WMe0R
fdeftz+pThh9kmJ2Lo2bI7NvCfB0ExVX6giixfILi9k+mkdzBPpIxyAy9A3O4j52VY8bt8Ul6c+B
dR0R+NVzvL8Itcw8mHKGSww3s82NMHjAxfL6UkCIpbw9GHJBSXPQHZ1AOOJDh+TPG72Sa1voBy5a
BHfLycibRtuV5VAY2DipHxt5McQAerUtoE9Slh3ZL1IjIDdxmowhEEfF6l6o4YhjlRK0Sc3Lys8t
K/QR4f5y9spvwdJupdFMOy5X7izi9uGLDzoBRiGOdbT6jfGcNAVfflYICjVbRdICA40tQ0MggyKw
UJysnxj6s5oA1Tj3AFLIZwyq322G32TkpENBvuFjWBmULb6MwEw3Kcc+c1/codGVyE0TlJTBK47e
GqeW3TOzK3E1xOZCrWgaNDCw0lW2XmB2D9nZspNj0Wbf7HRy4CzKYF4wCJW3RY4Gj02xB8E8otSb
UO0ro5vD6uNBeC27Csb2y3gEKC9zcIwbXaU1sa8C38mfuplLckF/O3U9bteqfmObM/lxwa9B9RKr
AcfhHlK5nvOyvgc6/AOIAmj5SOg0On5O8bN5Vh3EFwbK3ehzu2CLsukUIpayUxgt9FBAK85+kCMv
x/LH7CrIvGUFewbyVaf3M+fahPTDK+gHq8VZnIl5OBce9e99wnTZ6Nq+L0W+BdlD5I8dWsQhJzVr
ZBWEM5BsJ1BI0W7v0C1Dd6Lw+3P93UmXtfxLiPQqrF+upgT39FaHab9PHQwgMLQ1YGmAKv4ouC+J
PI/+z0DlAvEmdMnoB2Jk2CJD1kqyz3v+h3CDFQIyyGQYtIIO9XxUdAsw3FsU0oqX7GKCrNEbo/SU
C3+OCa8wYroOCEGhRTBJxzSGyKdd1d+hyxKDX/tOYw8ekWuz/7JJf2BjHE5yqt+uIRW+5XKnxi5T
YqneN0CzFkehAUvVWjmOKMBB9os1fj13a1skFjUc36ihn2woKWEmIrS3arLjbC3k2KLC8+JlaDcY
la9dcmWD5ycRb95cjdO5Uq+muhRYLCl8cHPhEeE1rqqAEt5KXrcQclIhlI7At5rfODlEsW6vauvu
+JU7Ck4up2wxtMoNwI8C72MdPO+9C5Ov1wZprwJjxh5CHLgFGijDKev/bnmeO0l6pnesAw8x0QpY
rR8Wdt6YZNMCIBEWA9RinitQkATo2o3CX4uVVXJqOUFfNhuZlltpzAjq48CXDEnWD95ssqn4WfYR
rHvxcFuDYpp8P3xT/c451lRr/VudTXZ7j61mHYbhcEEAXgfRHk4fbZ0UsDK2TxFmRMQgchm9gE6R
pywB3tSQu2/OJou56mfvNUifQqM/e1jWG23XmNtt17zeqgStSXvvnDPxGQyLiGcsh3X1N/52V2ZN
O4noK+oSWpzdduG1c6yLsZUFhe5JcmoouJczGx+Xn2QOlSICzsVfy9Siu8T70/bZg1vHk/oXLX6o
ATg0CGeJzSNgUB+eFI/lC/JFNBjgXLzMP42DXmRlZOXpEs9C3QKx+wU6xC62/9/v0VBpgQcwkudv
/PT/4YVK3+HJvWpXIGflHPm4bcZpohf/MsZoL9LtLGZgFdpGyqjDBJCdK69/aJEjM6mPlpLsYOj7
aCco7JJXL3eBcSkXfgvn16kUsRQ6SEomStA4wvPzVQo8czKCgJLznws0D49yjGE/VD/fpHnXxfYl
vx/q8E2Niv9k19JSLzV0jT8jhmWDhBCuYygA6YZowknYz5OPdLX5Bzi6MMLbJ4bVrlJxsHWBNeKo
LB2J1p69Mdpuod6sb7XrUW2qJkPMy9yhGFYYpL3CkXpC2rfbrupe9KoJAG4orgwAJW997FjQJJG5
+0LHXcY3oMdciYbG4pm2Y9xW1jMTH7LDs5LENYJY11RwdRrLn30xnf5svoLi30HwTU1qh2Ribv9C
SStq/SCtXPYW2vhqrTKEwV7iKTmBmL+2szJQUwTKwncFrhbj5NIhBGye7ZvtSiT7bzbhJhAVJ6Lh
J4ju6SE2v+lGFtyZMyhLTrdgahGsQlwrveSUW2fNCZY6xqbyYCYqlm+Jc2PYl/pIDRQhpxRMnRpT
8eTGq1T+WxG252LfWS4qB5OtujKnZyGhD//6XPA7ZiCIPaVNqCB24lQkxDVOwq5as/x4ecI+fIVP
u6DL/YGq8KCaIBVGX+lViYdc31p1SLgEyv4l31sFdcoFtJ5wFmpvVa5OkwXXSZL/bIPrXlKrO9YW
cthVUO4aR8NyHCAUNc2e43A4ngz6HKlKdLXwCA5F7ZNhEMjg1s1iQ/flE+ozG7Ghcv26NopiB0BC
DUFc5Qb3DRDIUQpp2lrSqJPg7VeQQCR0DIhwtW/iG9qScMoylmvDmWb73hUQaRsxiAWfcHNbrBn3
1MXMqGlCxu0XkWWDf+6oUwopQkY5zr8XHgDCV8dJh1mFtiNnZM92GqGkE7NEXq7a1ZNn2hbs/wbp
uNfwNBXtFAC9QCatb66S8a2A2crcDsFmhfvUgh4vOSdC2JOFlqTVSRORHpYrRq5w2bjP7u4Xy7Kl
XEkY7CEuRprNuACI3DNX5LAwF+fxlxGMlQPmL2IZl6hwWzaFbXnnM0DZBNWHDO40I5fuoEBi1GCX
2Coh0P+4DwpqKjqivcW+J3vJeiGNJ1WiY/yH1G8p6yri2vafQGrLmgd9bTQw0p3T3FyecfsO69Fp
kLgQlJ2pvpswmEcfa8VwjOHVvWWS5Nbse6nD635ZSoH26UXhubErDh77rdycubAqYyvyiwm3JFC+
rp5OllbPdUsVNuGx9QE/MVdvqOohnBo2G7BLoCb24bmZk1qo/1zumOr7KRQwESWb1sphnP96LDN1
CNWgyr+Zjn50QsvF4AvwDj2+72ub7eeHYGJoKIRlvP2/QECkloOBbQgqebFueUGgzAd0yaEAXnrd
w2Mqezuub8qQM/YAGuG6zCbux/tmL6fUw2TCUjpEJQ6iQCRJwxxjF88dAfID1KHgx9ZjM9Ah5tGJ
Tx/ZvRYy+prTnA5uSNnjx9+SWCYVww4XqVWmp7JkeIvijMch+9HK6k05XSRfSEkxCBl/tJAIeZfT
SonzWz0lPCMhCFGz9lMQFxr1wo3aXyXPiHN0j+ZxbcZVJbNHRxZaiGepOIA+P0p1heZeVM8US0+7
my8dto2OMpGuKCYKB3zdvZLPDlhP4kwHAt1jvoN7+a3Bmp9xawLyi7Bni/cKXF7MgQIYIsUxdKHy
O2a8h+WanCQeI1Yjl3EpETJxRhVOT/mf7956JdJuptqtp6MxnvsmokQEvEEO5AIRlJbtHKLn9JJl
WCEf2+IFLQpEwSFs34onxZBft1dlkBqMFOQsQQfXTLI8kzUr18IyiEt4eYYX3PaNSN7ksYdXiO8f
mn/9AS6rN6VcdwHNG+jTijrmo9j0f38RDgs5znjm+1O+BhmwyGBYR1x20EqoZwH/hv39tdiQ/8wl
gIqNj6Qo7cRfdk5BsKGLXI2nvR/fZYfvMmyrcyM4B/1qmAWbDEFJiX+A0ZrY1tVLo4jgdO0Mpvc2
efIpglhrOKEXZImMYzOTgFnXwH3fe7zB8RJ4eNxu1bgN3/Bn5IqWcAoXLv0Al1wL1yWv9XFBy1xx
MY/fpMJPNUj8AxtNJR8vw4V1uaKvGURBsnas0ruk0qb8ZjM6TFlPwMdo7jWCajoGoar3d/mCFMRX
GfeE9UDv06hshj2yspmHIZPQAinopNMEhIVB7GpDoVVcLcZo5e++GayscidwDaK/61l2O2J7yFHh
2lsPSVyU2jL30NYyHMLVKQwZ8rO3McDpMeLwlXSUapr30khEOZEFGQWanBeMp5gpVsaeCHISjV66
P4ASyKcFLubsTL5s0OnS0ygtQndZkbenRuyvOHhH/Zhopv2pJbHghO3pH77maU+om9cfgOfWI/37
G6sjdoT4Im0x18FE3fIbq79NtibhQF+vk8hHo6wm+x/KeE19w9/W8nkzDfl0lpo8G6yk/FConaCY
XfvddgOVcD00r0l5iYzf/z4GrsKfwW16i3ASXGy49R82PW3nwtlOGvlY6/RGt3BYrHpplK7TesHJ
vBljK5q4OijhrDMh55siSggz3YvMFu5SfBWtcnfZz3DGW4JSCYsPUZ9IatDOdXfU1P8SZdlGe8fi
hWX7GS7zTvdbz7UJIXefySB8mniRtFG2uocZbN7p8CNKLa6Z2XR6UEJAblyCa/Psr+kJin2oAEHm
ysvEC6EvJ4jkum0D2HekpIsOjjCrQqjw4CqXmOmj3hr7r2bSi47Ge2eGK669YAgzN3TFhuNTl5WA
3Rh8Z/hJT2K2uCZLRV2o6T+BBi94zSAGnQlLiaH2EgwhcbEuUPhlBvW6NV39/EqMF8r3t10hHmmv
dWVsM7kZ8T6TX9RymeENCaxpAT6/yNwwPv3iKrvQ1CURw6YSS/Hz/r1WbVXJfVtNOSVG+p9+YRqK
fIssMxPJKzkVyUIT1kTEcA1N6CZVvepPbUvZ1Ruigt52p2YrDEkJP/cyR0UIx1SyCKDCStnX1ELJ
aH0lJuVMd7X2yTw/CzbDKu8gJC6rXtrq1ezuTbSTZYxUDvfo2mJY9xo3ksppWNmibw43gWIu2o+M
4lIGURwF4AVOn4cyJW0g92/KJarxtmXjfup1VD0zjMQkGZ/CqlI4EmK2gXIDSLa5GMoZt8FTF9Oa
ptKbgPgpuQ5ihFsrxX1obIsUC8zo6C9ZdES0FLQu6b7drexQip+vS1XlEmxRcaCn+zabWqIZ+qDA
stt9vixEdwCJJMRwJksFqIhSBdh+s7cjNJG+0/VhkC9IQC/kYhbEwHfg4QQ+EeI7AB4rtGsMYJBb
6INxRiQx4w4uytNLsI63V/NjI8eBSxw8IG6xQtHEthE2VaY6j4C90xPnjqxmAUYNU6E8EOmaKfp9
TfOSz143t/cJX/YQGSwS7uo6r6JskkqzpLJR+UyN6pd3MP9sJxhXAWYamLuI6p5uvjxlyv6hTtaE
09MPSSFvo7qF2Up2kQAAibzBdZ+sqdOLieqxvE5jzzO4ritCsRo9Zch/NKG193oAlJF9Nrq3dNa1
IixnUVyL/P0mOnK5hiS5TQRpN7iCsedpyprw6VdY4QME+WVaYLSElsC8wm4Asxpi2u66IeuCgw99
XAYbAZR3/2yk53DuQaQlBhK1ddmGSpMF5MNeUYKhK3+0QPLuR4UjeSL7sxBGZ7VOR64iQlz0aSZp
ENWpt7JGEBuZDZrwMFe2yh0awkXIAAFFObgtiZo1SmCmJoT1EEXy7/5Fkf0MrN8hwzqeS8n84Cdf
5uM5prCetBelmr2ne3ox9kwF0mheTlsd2wFqEqEohAQT87jMDaguflFBwDAOlhq20VBRuFFZWyJU
o36zhJJKwgYf4CiUHaisGUlv/yJhQTneipSEZZ5H1rmuWbWUCn2j+7Mk+cs3tRkm3XiqPYHRxlib
jHsQsTuh229AfJ9IxfM4vLcbKkynVp99rAA31c4EqHd9Ap9sr95nV+45Egf4+iVlxs+a3qR9yOe7
Ukx0qZ3gNKMTRPcqeRzmi99836QiUGJPEf6lqYs01mWw2YRcm94sehv3zUvqsyQ1OZTwc0jPWMo4
339TIYI4R8N1G87bPnDpgLAf16hEcI6u9cvM8hWIUkDc9kZDWUDhjcN8PngrZeAsiHrdHssRwk55
xn1YBJZpmblcDk9UGreZu6VPKs7Hfz+lYFJ5BqYvwUMOaqeG0xuPULWxSz25OQZegYPaixTBmjZZ
E7elhXmFepplXZPxZ6FSl8/vvPzkkrwstK1EtDWjnlmb3mfoJidV5fIzNszK3kN2M46QvTkS92uz
vvyexYnMu2zJElm/Bp6YhNHvYTZ6wV/cOMlRj6+5IhQHEtrJRQ3VxQDyYsfYa4jzK/E0e3O2sqJa
XqzYMDK+bH5kV/ShT2j8hHJsjSv9JoDzts9H37E7whFB3tI6bcPTEGnImXV/rgHXM+6U0tOV+AbW
Edh+ANDBcTeXQAE9EHRuIotNkoNl6hsodYEhMzojU9zkp6FEecvZ64hMFxI2AixxCnn15tOlPOLQ
GAORl8Zk5TriB8UFPLr79PlW5a/gt3+6P9KIrbA7nzqyVJ+nZiZj0R6iOfF2eFP4Rz/WXBbm87eI
kyArfzJ3AdtO/Irzw30m4B7YbbQ9G8T7d2dbFkGFV1BvM5CGYZGitprmSzIz9PzXGUV5A1FWbeg3
8HbXP2VB9sjuQ9c/hXQn4sGSBL5t5TnuTXQzp7+foQVNDRZaSPB7WD7r+AbdbcFfzyugXD49/r2G
hY4Z9i4zTxPziumLC41niI/U5X4D4WoT7cVoDufNWYdSkkaW5KiwD9Asl+0myXjaY9i5UDy7mLJ4
/JB9bx52TIGL8/L1M55oE4lDgV++yfzDSMG9SubRXtTMz2y47KsLmH3zkski/5b0pmFMQSfeyEbB
H3oUSV3vn5pDlKJYqvNM8lhsYB0IMcf4K6ahG/wqVnglBpteae1859bDGwogw72ICxLOeYO/k5Pt
91jUa7JEVV4erIU0c25+0Y3DoBSnCPDsT8YivUjhhL9FtoPoIiLHjveJ8o49rTTWWlfay8w2VF+6
hpHHlhaFcW8rYO/5rUszRJ8cfJcw340Fs6DosVGzkDwJMcuhQrjk/hNDjcbt2LS9B+ha/IUkJQyD
uPYoslwGSopAgdyUo3hEjL8FH419VjM9nqb85OU2EC1V7Seb4bCXH5MT6eWGICHljNBE34CGDbNY
ASrIXIuPDswNu4YnVfHIvXdp6beGPc8dIifH7K8KAA2/S5RiL3351V1djlvcMb0UaygTS0q5Y31X
xzdj6M+Lw7A9lNfQSwBJfxKk8dKcE9IcfR8jg3m6b7gvD348azclyVu0mfn2GcWI6sf7JuJ2XeqD
Xts7eW5/rb3j9I1AL+XZjJmltBRZOP0AQGP6rjJZTlOX02N/UTl8V6MhEt01UECEYWmJsmFEchsd
dKd0PHMJL4fQ/j9JgXfX1oZ2/d9VHfsqmu0SZvMA523XbIiIOo+K9eloG+AS7eHFekknUbgF8zd6
2YkVLqCjP7cIySYIqPIXO+jHaw5dFEy6mRvfGpUuvpteLtX0m6VAuFZWhBhY4WsUtl5g/w6W7ynj
q6su7XzaRpwVUr+TeZMwyVaQn7t+34sOpqI53Yt9C4ZWJePxNCTTZRDNIHXziWdHTJSjfcfDaVmc
5nVO6+qNkp+nsEiDGtP0lw1c3xhUKJVnOKHaNOA64jR7kuMH6390rlYJD8UwZ0FE6Zwxxxzzb5Lf
Y5ci1tiXw0idgxI2vqCKTQFZaIVCquYXJ32NRw9kihO85ZM8/BV8S0y8bqwbooKXA9xuYtk8xA1N
jtP6PCuJ2mwNBpC/Ts2J+Z7TUTmR74TnAlnT89ALkESi3KhxfLJ8P0Wv6n68bLCNtpe56Db7DHm5
wwlppHN/vt6KXXZVsaPJIAoGXh7imL1EfvGnBPaLlRrrPgLEt3TzQWWia/hDGf5j3c6q2DXbWLqt
o5PiTfUinJiFfPCeypstkug7AITUQBDJcoG+MDV+j/L5mTa3xUvby0TDSlcTqjwiXqJNNp/+h4a6
ubdS2GdSHz/G5mpKFiLRWa7eFoPqLWtaI4ZNb2uWOsdUSW8/+yh5dV76NmLkRMv1aNfGGRDgLkZf
zUK3SDjER5nKlKVKHVZPP7SMSoTgq0WaYHnTxfav/ts9Mfo9QA6btZDaefXrbLnW5Nmlsqi7yfQ+
4SKVwpAYUlnj9d8HmV9ofxBTgYAhlymWHoruvhCGJ1UZ8XNAI0wi03CB77gVQaRCt+yIdjexw5/h
4d0UtHOTe+/FIilEtKNRpQ1oFoXuWV4rgASrQghDQG0QYxBo+JlxbL4AnSYhZtG3NnUQnSyHRA48
bfZogi88/Kt6Bh3O7sEcN0q8BAZxrrOZgLoC/Af2k5kuPAMH9c+rWgP9ApC+I3mNlyUVp+ZYJksW
3dfrqO/RFn2oTUUjvhsaxuwvwmAylUb8Z4NGux4NBEyKyBpDAPDl9U4DIj3Ao9FiMc1apImOaLBi
T8PNfqX1zku+BwfB2G3AS9fOWByuggyWmgxqxzr0ADnQBOne41YewyyZjz/5BmcGzyfg39PfBf+B
sbd3I1aHpPA2kcohk6Xf7UVanajn63c1YeC/LX0OKnMsiJ5hjh9H7tq1IIcqJZr8dE39LbLy7wvU
1Gp7EOU6auWbGgAmgBRkWOuscPA5wFJ0Dq43YCErOczsm/N6nZU9X3CBe6ECf6UXyr2hXx5I/knm
WRdikrFiw67Y3fjYyPIHg249sbdVxKQBhyqcm+BkBjFBv40BD+MjOcIyuJPvfeOx5illHXRO+yWv
H1RJW/vkuJT7D1zbqe4DdvuXs6aVmh5lvnW9mveGqnVPP2bKNCXf5h6JKKGli1Y6+DdAabfg57vv
Nz7AHtDClPaJhhad7R7TYxtVP4elNAYwFDKidKZVreJqrENir9DP19YNpu9AXdfX1I8rl3MIWmKe
7g1mPlV1f/RiRMN/0ettS9ywsYFtaUI1ZYh0CUuuYHDLJ8L8MghuK4dlaN5P8sIGlhbLupa9RLTQ
OK++Lps9VKxN2WUywVyae6K1xyzlx4egLJz5gWvnIofK9gcHWVHoV8qokTDF6Uqd+HWNJi1FLgjP
rLiCk+n9Kyb9EE8c51MzV3msqKkThU78r1+05+KQDytNOA0we+zIqd81UP/lmvV+JfmMSdlxO7q1
y7auzK5nXu/zRh6IreDt/N+wfR2nQO/flZATZxIqveNlnlAujg9+mOtMUPjrVQl8ZbcBnbnV6WE8
dT/VAb5ejYiYknP/4+j3yffoP5OjJyyFGWshlKwM6FaIULHr1eQ95tx2y8OjNd2tmMDEjaK/83U+
vjstoQyIgz3gn2FH4J2t6iraFhr3nI7VuqORrhz+L2XCt2cv/P98/bczF8TZvaPDUcFlcAU/mUJ4
7WsQFwhnY4gDY2coTwTj8HunLZOrPkeYO8djkgs9gCc3SSpCJFMzh1c87HExN5ExG8i3nQRR/cCR
3FJbPDl4vT2Ac9pEbQNdeYcN2ykBe7oBh/nZXFwe7UJVso9g4p340AtyzejQm99eAwggwzcrkpo8
hxmZX9Ffs8Ii+rPOfqTYBGxu5axv8FoV5u0OErGta39IIDH5HkMCwTSxSJccNilEk9pYc8hqevsL
m5rt81KjYi3RUK4Wt/BTJzLw+9nS3y/qExjNmI31gaW8c4h+mlhxiCx1KZ+wpqxWyCcgHvnVyY0H
oUO1a1EaPmBgnvZeYlWlskn5wyq151JTNIA4C7Vw+frTp4s8RdrFxb3U3g8Ish7I+KFDEkTlIwLq
qjLg2OSm0kPuOXnUDKH/gA3T+wq208M7SukxwlZjO0D7kYTMuYX/4c+eTF+Ktrmz2meYr6VxRKn9
6oz9TtRXZvvLP/nwBA5/qBLgESKOSwPViaCP6tVzaRChWpFlHA69f0gwd3z83yE9iL5wzKrYWGI8
iQAO/fCwm83E6n6Nttb1+oZ8hgBJWH3uX7NwTYbaoKrTgosoJcvsUkFZbjImPv/SqePCiMiL/465
v/yBwMmqDTqXZpOAulLl0IEmGrmedfBf6KtYyxFgbaIT4dYmM3l9WLrr3AkxsRMCkD+QCzRAB7ss
Xc1+FV7W0C6Gxc6EkHSIRj8e7+77tmGGGVXNuRfBluCACOb1HdeYXlUX93vKvGt2KkRfgeHaU/Hj
i2eCye5skNtT5MujSeg8wzkYj9HPqDxIgaGhTj52zXL85PpJCitEqLv0nRnAzVoZmK8fiZ5ZsiYs
y20pFktKvxBR4g3OQQyAdo5+3Lv/5ilOXULh6wHIY1A7WJB8mmxXW86dlca1iJtuW79YPi6JT5MI
tFBvpuHvcUyprKAhpIoD9xtnx8zAElrRwxfoXz51ZD9rMQ5etvemobl5gNXfC2J4HNEzgZGXYrLg
wCwIk8QVrfZoc+yAl5B6DR85/7ppk/sF2q2tzdoS0/Ylf9OlRru07rwmkQx8vYACowkQ1gynon+W
Udqr6NhsAYjew0xZI6iyJ/OBsu4FiMObr8ylqVhLcFhfZNsPYyyATHHvm0uewVGQv4GfEWzukV+Q
V+YDcNgPvJg4Hhj3uVRVbF5P8ZF+YUfaDedPH5ZvD3AxZhr6YZ+qsdOQS7OjLdbK0vBxvni4SjWc
K3bUQMaHHVM3R8y5RyaGG5pPhMzFObqn2lVCvvOqN8O25eaDWw2MKPOKgtvlj9ozw+Ol5cCLb8SV
+YN/xVFUjYnCQpOJ4WGpEbPLE/7fHDfimoej8mYXOUaGq9cll000aAJbrO2waQsFLRhdb3ssmeof
4uGgCGF1DSGB8d8vaN2zJtV9+bTbYix6VP275XNrO1PGycavQlkIanYw+uzrS4yUkLOdzOI1Vy9q
tE8+xMYYQI3LFdxm4EcGi4wfKshKHtU2HyTJp8YGDjj17atZ/RYYOmrB/D02UyRraVVptFYQmSNF
GVwu+NmPcvMxe78jx8u5bGnTTwJyJqHhpdn2VG/hEZZxqJ7xMnjRkAUwpS3VJUBpHczB7QjqQ7GO
W2Y6STBOCMKEkwbvny+RNpBmW3RgFB40lKX5SBiSN0+GlQL2xlauoje9KV1cZfe6+i4DkCGutu0V
gcThiQBlXwLyesW7kF6lNFArXTSZGLcWG5TbZr2oO/nu84lJft+viejFnmdBLs6spzESiuiakYZW
3eQ6i0Sn2LINjZaPn5Bvn5WSA6TSFbwAIeOHbaVGKzIQinDglovv4pPNL1vaY0v/ynNuBsVtvx3g
UGa8cuAMahceOwLASAFKwvYUfxPMccwmKR4wknoYhab6V3U88IrQNFwKZ2svyEoMq7CBSsurflBI
iEig+l86Yac1Lt5Tkyqmz9bh1X8KslYvHIBIV2/IdQ0xh6topWAchZ8lD/5tuLnr7t28AJ14LZTT
U1byZdR7eNtQhhkrYlZsHr14UFrhEh04vdry6DUjGeeA3AEwAHSSjqvfDFSIgrRmyi/Q4K0u1Phz
jmLqVGWxK/74EWJ+ke+dZ6sqMsIOvfQNUF4Fb53eNrCK8z6Y1ptaR8RiTnRKlbvLOA4cabO2aNTQ
rqg7+PMG5PdvHJdtgtbAtOyAXFM13gn7wD/C/OwnaVVsbJwJnDsP7DrjKFZh9JlpFBSywFXR24Qm
ttVwim9tnJKGLbY8ol6aN39F+PbDuLLd7A7oZCGFO4VCOiVUuFImvUc0RGNco7AMB+iLeUFpUA87
ledCiYX25I0xrxuPJYxLow359RJmXEWRM6rbfq2qj89y0Zl8eMRaV8b2RJfwLxOgkcGnYdLQ8Xur
O8tjCUr+RT+xmdXrjKcHZBPO/LyYr5vzyZ8DJx0zOfTOwqBq9M8H8IPxKXFJLVPvaLkHiLqBinFQ
WPrhN5CIUiIvcC0H0ycA9yQYIaR1f/g5KyY7oCNpgNHfEsznzQ8y/DIyaipJ1Il2xrUDhfxG0oOQ
SMycW++kU41XsJhmaQNzBdfJvMNmSzUm1l+INNkot1eNiVDcztMPFDjjx/9ERSoOLtax7v2qMOJ3
T29t/9ckNYivuwL4dNwU/CLOCPKyPBKjrR3jdKcGdWEJkUiLvDX7TNq6EFT1oOhXnq/ZZkRCfqkI
2Hn8bQ0GaMmZ+uFfVIJNWQmSrj7k4IB2Fldoh2Zd2ayNLTZm1938yGfGyelZV0OOVWdH2RDylOXe
HTx9ulFHwtFapIIuGgUulHkbYxbfK4upKM4xR8DkQUZwuuJLiqhLhBIOsKymOU7/1MODv2lq/uRW
oycVZui4/t9Z7bsBDodsffkRRAsoOJERP05gT80k+D9yCfSY3/lvbC7yguwnNM9oKrHGjmf2VwHb
2Vpv6/ls5YfvcnkwkSN571qCNEo3eE1xXmyn94Fr9N3xEGgma2b3l1HG+gOf0TNprIkBtafqCm7O
LXnMj99EqV30qvce6JPlqFO1xmN+sLHl6xde0lRhiJfK/lrsLeeiq8srESqODEnwaGGo8mfuC1/7
j1WFX32Cp9vB1HzlWk0GJ7Un+VQWJP/P8DNvHfcjJekvpebLBELnxgctrmPrgGdTpBwlNUbYq2by
NSjMJckuYh7ztYw4yEnu3QK8LSJDGKnBoSdtC2Q4jlxxlguVepdD2w83XkJrLqPZ9EC2+B7qU/i5
/XPx4pI+R35GYVeGplUk6ylGcS4zQquwCn3X+V+N3DBfVcT8EXAUeHJ7EENXHaYA/OMLSge6VSrn
4mU9BGPsiRuPPQjUL+wHpgjFUoPo5rjkDVWSoEDxq4U947+qT3X87sYg+BDNmfVQ4lBbTBE/Lsl0
UFid0F+C7p/gmnH6K0q01CsoYqj16FgvMdyP8c4yf1ngQBiUQs+ROU0fSPB5/HuH/Ou5hZc/XBun
4tp6yiH7aQlWJ/LTiH1d4H/eGaOOQDQ4dJKl2DDCrccpVTheHp88w1gf7rhJBcHDL58z6OZgHQZw
9lWTrKGpDXOySYQIMqKwa7mYJk4o9Fk/gC1qit2OjNiR5Uh+7yfJ66SGycY3eNmoPReCZsGHrxQU
f8LS9G2sM6f3MO9wCy2WkkM/DAINkcCwpRSxoiZtnai//gglRo9+8xhtE4AI7wCTbYFD1Jw+ZU2z
Xa108KxLWSJzAS3/zAdttdXeZzlg32PFaTALJ8Rr9TAI0KxLbQ5r6Hp6kmhmS8R4zG3uw9str+63
fMH+sizHLGxh0b+XsoVp3Wbi8wSvn7MpeNR9EthJJaXvgvJdM0zeM++xEDJQfbb2WnMJigg4bmQ8
8lDEOLSWjEDAAzbK6d5vbZmQO2SA/Hy/vHyrOPLNoG0Dj3MRFt3HOcFwJpZorgLsTrJzOIn2oKFS
5xZVfzJnZ6x+PQl+6aqqat1O5gN1SbnukV2/3LM1WIfLTdiampT4p7/QRbmiifBXs+7tssWQVxl7
eR4MT7mc4ZlefAVXGEMild9HyuFIQ58QLW8Rgxv0Y+RuanBn926Hm0QfYmcCUvpqYcl35c9slSAO
+P4Ynkmb3pI7rtYNlCCXXMi4wylEaTszf78V35zHR8c5STSQlgXwzavr3f1bZLs/ZgFTh+5ceDpj
VhFIhPencdGhmCxSRvaJTYDztkL6CGDZyhJcvcJrKowTlKRfafqqCZsCbRMX6MXsxOfFsyOPJqzK
ydvMsRA/7aZ2f0jr73tlhKsHmyvMrWVAppkHPL034NjPRjUjgdkU0KXvb7NktNwM4y++anegjIBa
FUTuhj0dSctGlqWX9A0gsjctWMkTnb0yyY5FdWWyonIvWSnBd/4TFRhUq1NY2rsbKEdN7BBI5Hm/
zFc+IMqSV5x2adzJ2lOtXxMjQj4hGKjD9Sez7lDEbuEZhCz/Ju7tOoCCkQJ4g73DMGLhDTzbA0i2
1K9V19oRCBRTykG8E7887XPIYGaq9zJML61LDSs8cs+/hBDuNddSEF5VyshT/7Qc9aCXCJbyyHQN
Yw7C2NQurEw9+I8Gsc/M1ioghaTCH6fPs97u3d0oAx73MWLYdnfgE/h16Tl/mm/n1L/OaLQRyr2d
7ah2yzHTCg1Aq6XfcR/PSs3xA5b4k3+8kjt9XV84BduOAk63T13WvlrmJjoHKmoST1hVsUU4rdw1
zPR1Pe6j5Ifo5Ci+jCxodCIWWitN1Tcey7rQZcQTtasLvKJfugvXANxYBFUwsr6HM2XRs0ei+n2c
eFWAgry5jaf7nW3A7S0FqP5umOMCLXdaWK1br+JpJtuswfT0+jjT4geKF66a2OsBQQ8IbruUIYFf
+0tlLvTndk+TIsNuaCC7d9D+6DokV/L0vTJdhXnAboCPz8FuBaHpisWXZL3oND5Zq8sOKvTyHfwR
4pM2KgQon/4L06ZjWUfsFwn7pR/lyiG3dRRJqdHx7TALyzMxWrQHeNw4Nox3GWfrK6n+63yDFiHs
f16BuejR8bLBliSOCTBuqzDg5m7TAKtSr69PMhPy29rpdO8mZQFOYeldveE4SugwNT+wIEfF1dHy
ZTsgO4StLqzcdrDsnwyKZO+3aaVMoujZEJi6aPc1lS8zVZDiK4V1Pha+dAqWfo0StRdYUnHUqYyb
GIX9x/gmse9ZoqRLXh+Fy4HC9re/GScxBWYGtEk5rkHuqw3W2iXXX3kkl2bU34OWMLEaRsxa57gT
Za4W3RGCXYEnTNPo04FQmMH+FPBd5TnFVkCln/YLuGz2diNnkZNZXz8S8gp11xJQz8XoltePHmzg
KyiuRacDTvVaUHau8kLsh6lIBPlY8+EXFBEf5u/fbdnFW+lBHxWj8E458UDckcDrz+qfyVG7xsdf
LJH/jgx+x2DgIz1QyFBU5nE+UmMXZOIKJgg3Oi9REEb27CwElPJj6VxEnntGGbFs81n6cU5Taoxr
AtIfN5aoZjKW7rVfouko3XC74Xq0uc47M50fZJu4BptHLcXhrSSJc4enLcLqSvB9I1AlDxtFbK4L
RPrIsCXCQLTkqEp4QX41JBRE1S7u/iuw57WGoFD6RQUsqUI+SLnODVhsnP8NWdmaiQDzyA+EzRvk
CtExUJyA5sgP/mAtxNQpVZRXnp+c5jM378tBQi+UqgJ9THv2b8MYelTImgEa6+o6/8yRKjIEW0Wk
AqUrf0Xlmq9p+BRv1Qudj7QxBE771jrxuJm/8V3oOo+bBdKVyj8L4nEsisTtmyp+QUfv9GkkeZ1l
TUhmc5VPbdOeE2r4RxJU3PJ4u/xu+D5ZqQB8a5PTywgNYHbqvIGXr/VASABEqAZ7+ffwh7JGESGP
kqlHSmlZ2/YGNoKB502yHiOpdS0BLMPL/VCB+Qn8jDameQUrxAdDCJbYi35phE1OHXW48891kYb3
ib18h9gJqPJ3CBsAToEnB8FTFSY0hYevyhDp97tNtUsowJpXNLaTCaLiBcl2Kfq4bMN/5ZEkW/wD
h2nl0YMeQ6Rsp6HV4iO6Ewsh54VdVI5wSdcEyEIHp98lVHKS9oRq7YR5E9fsPzSOQ6MetjRCfPw/
/2YNTQ5kJ2FjSzQ1Z4NXT5K4srdyjgw+kCSOekm4quxtLfDLLwavWWgBTNypkXR0y7UHgVgGsYsM
4HnJwwNfv3XYwLgKk5xHnZZA/ygaTmeftX+hu4pN3Ccfcnw02Ulp4sMDQOkAqZmvUs4wPZknMnhd
qKSl+KUeW/q/lDQ5neK+JNVOHk8b5LthNUG5R+DQpO8Dhw42CxKhbuwCZ59zjoZewXhfKJp82Dfb
WNhEXTORDHqF+h4GhVVVhm5Zuhx56do0gOlsOzhVum0SNXeCDWHcpTejTNpbzD5dDtrjJzJrCMFg
QjVpE5RcRUPW+y2ZOKb49Aci+YITuio+A2FNn6PjVrOaEAZugDL1kCajusGmd+LdM1T33oB8///y
KZNR8Q1qrmDl9hcgJVpGTyjZLYSvC8dy/G1EOadzaMFs3sPQF6eGyzR0x4IjjQGsgmSN8oJzOju2
XA99fa3Cu1nC6Rx7OZVZmA9SK0KuSmMSZtRVrThEFwkeS2mEtlF8f5tjaWvHPdWt354Kq2m2WQHj
bRQ8HwXIe1SnSKyXI7ZEqvVzQBcWjuojCTVMap8dk/oBQ1LE95AYqLb4i3nD5h0kGG7JVAJgtPES
mfRntZOk0mcZKdeMH3czY5KrT3i0AgZTkN/P5jFKDLZa9AjyZTiFOpk39zD3KqfygQX2RgbS7GsE
qT3N0wyJ5zGOMb+WXRAPTzQJOElNaBtycWIUl7cP9UN2pVC1TtVDC/yU0xZzL9NzuUM2vTIH2f0o
euYw5Rf2neDji3caQhppvsvwV2jcbGN4NYLcvbQaMaRta15kl8g6RjIKsGf7f/rYwBnQqn92OSIW
3Xj2MZaN3fpi1ay+Zxh7pnmKkLQYCX0irbHQw/AzsU1GI6pEuxI9DkUiHQdv0FXnoxcuzlH6w3zo
SQRUPrgb2hwCM9iSpBBWUxQsfRQI7AceYSM19qz6mcCAg9wgplEUUv+qKYsw2IBRmFuMoGWvL59G
I15v5Wpjma5OYj0JtaMrBEntgE9Qi9l2QAQXSVdkWp5xLNwO9JQcU8ZJbIR3vSo7VqniYNi0xe6P
lf3I32jtq07z95hWCs0PD7MDLVnoi1zixDf0u7vC2znhJCTXbciXYVFsNJyHih9+iFMFHB1ZX4xi
FDB1j0+a74pgTuSaJIevi0M6vuq1+acq0ENBtxo/NiCvPvJ9P/t4wRZA/DiJEganCPBSRPMfmIAe
gHq70ohLWbVbqtt9enk3Xjn16JKPNC6pxDa4ITEEMECHi8zJcDIovSbijdRHS8s+IfpYDnYUkTSy
jF0oaxIQkbMx28Bh9Uk5La9kjB7RTDYEB9tBzybtufzRPoeZw2y9a3QYgPnWmBKMXlKKzsBVkeKF
E1uuuYvs+fIPoF4MZPE+A8dLSFY7NwZjIdoDV+h+/4eCi/3AnAwGfbXZlX2/IXOavi0pdTxxPcJV
4KdexKyNp9KDpWOrXLtxunHpWK/tNnhKPjHge3/r+5gN1bPp5+fHmsTfIURkFlHT34z523MEVfiG
ys+qpBYOkeaRdwJv7KRmukPfdRlxoo/KRdf3iCQ0DQmpoZpGFlKCJQky3905kgV/e8YZ9Qx5bRiw
WgZxkY2pq+NZaj5KB06cRgzpXRCG4geIwiKcR6z1mg5w08f5ddoe0vNUh06lFDqgxIgdExkgoZXc
TUlayhZgYtqQzeklt572t67IN7hzgdeqgTJnqzIUHcdSJqhYErWKE5NpodQMRI2pN1VfzUSav0bB
DCVtKScaPf4Oy8r8tYuCZ7VDP/N6d1SbhY0TdxD1xEV+nNQ/WMAP3azdXKHQkTQxaP/1sWIZZfD3
OeXyobUZb1PmBOjC9AEPazDgdIJkVWx1XuVFOv8drATffUfyubO3qFhTaqBwsplDHHfJ1yoNRzOy
1ghCmrqoZ/uWgMT8eVOpxiRtwm18ssO4zNmPgIUrHxKjvkMkMB53gurThbIzTusknsLz4Tvf5osN
77BGQLmHC2rxc1ueZOXU49oPlstQVkaj2fowCLoifhjJ5LC/9vNH2oh0HtXN/K+G3v+exLaSCOSh
WtXItzU0JClxVhFONqq0KjwaPtTsm3liRV8yXIXlmpSvw3WvvfP21R8o6KdKL23iXdsPEmeY5ITc
WKSj2KrxOhntsR0GiZlWTxo0mhgymaJJi4A6/KicxWV8Aq2garBivSxeGlHGhOq2gpx8HGIvW/CP
ePSyhBKKNJqt8vU3YsbRRZ0xZxZvXrPNvJOnp60qqQRd1KmcK5EyFyt8cSoH4e1MCnHQLDcwUNLq
HkBet2eq/J9ULQiypg0s0yBIiseycUq5+k/QCO8TyQ9m2fYvauTx9cDT3bVO+ZgEpUvgQrXhZeJv
R6rU2mJTiYoGLzpJmYWzNE1sjNSCeQsscfCUxsxhlI8FxY3+Lu8O+Q7IlFIvRYHQBXefcV/RAYga
oxk8hZ5yBGePhtGYecibrDUsEcM/KUN2nZLBdwIMVxT6OogzSwlNWKZGUF37V3wFGOeBa5kkj+vD
csXF9TmGnhqgWTK3wZqUuc18sKHiiZKys1TfjKohH5VtlqvjuUMfwHng8jAL22Wu2l+VXxK2p6dk
SaubSMfeK73rZfynou4XpVjRDwnUd0EcAzcfrPGnI6DSNZ3r8iv8oM+YtMV35JF14RWjBQIVaTYE
tac0WxXgtSEJLNueHHygoO5JIFfitilX5NWY6Bgf0Lfr7m/A0F9OR+9Mdy87TdblXj1HsjCc057R
gfVZz6SVOU/Y5QFZN/uEOzfxswTvpMymCY7KxfZ4IX2krZVtC4CgluH4G+mLPBcJCt5f7V31oJh9
BradIGnZZoG/uXQexF9z844iz0Sq+ei4b3DZjm5msfrzzyuIf02uXznzQahRDUkfFHyQ6zCZOT5b
bz8OyJ9Ij6TvmJpEcHVwXs213VJ05oMLgPDSE+kIUwVTWZnINL9152ANGM0XcAS5rlv0jIyii6HU
Uw+j1N0uVTrxQAIryg3YRnbnNPMNMXUlUGNeXefUyk96ail63lehj/HIC1EEIQ3iZePGnBEoEHRj
i7uGgzL/nbK9lxdr+HbH+fGz0AF6Dvyxa60qGrhHbn/nsct1frv8n+ytEewzEQEYzD3C6+sGkELy
cGKRePmyv7sMH/k90LRCOh99c09kVyzY8zdv2q5sUCC0Zo2b9/kPjwiUMg7arGGL/Y2roDV55aQA
OJpAMQ1lAz/6jtOVKUznWVNlwhBA2BrBiHbo7GQT23ZvwMXmfTidadGe9ovAD4Qde6jil1ZAFl5+
2K/n1fK7zwX3WS2kmmJ7Hky5JoY0nV8I9Dci3TTbaPcbxm2rSyyia7gjr0WtuNKHyaaUFUA9hjhL
Jg66JMejLoTzrFcmJDWHPfPcy31wrzn2ejrZk3aEP7lpiLYmPR37pfjVRipLo/wZXmahTTN1KUlq
SyMcPfXnmOq0FPXlZx51cLk17js7iHb9eD6SbSY+e31VYNWKoSK8C7Mb1WUZ52VRao9hlPyRSNVH
yz0zBrCXBDDGvGkOzpqWUxuWl/17ykV5fDVze9Tj2yMEiCLaHLUWA0modfkL8x1u5wp+NF6Kd0FM
je5v1jMdSeZ7zFrp+Cp1I/b2TKGT+kJOS8w4qLZx1DNRr3Lilf43nvthEbonH12BXF5Lp1jWg8G8
KcoAPzoy42uPZDznz3YGntIwMjL99RadclwOJHq5N0AsvYcSBserM0xD7hXDbuyKgO3ahPSZp5ZS
SVWzIOxdrLPxHNZ+j8LW7sVEVf4KHVPWEi0kXr4xMICyPjVYQpRY1WXGKQyFLpf/MPc54vWFUQWY
OXYp6jEuIIJwb2Cena9s40twZV1lt1oWcOi4n+KeczTY+vLgYPzAUxb80eaWnjQ2VvQZciidWQkT
eM5JZJVOb93zPj7G0HYa99qEjuLKxH6YET6U5dq4r316sTWLB5HBIP8W5hODQppA/a0dqGu1H/Y7
bk1FQcVTTqJ6xvWi4akzlTTfBsRxYh8TtIcqBplyiY6d90PHvKP14oGAUppDH5NxmVGm9xf98pM2
KJTOwvhJCrflN+JaPK3uI61sQTjQIYyVtf4pTt0f0RcPSVNhe+10FYQVhGRWu9lepMJJnPCjMssW
M8C3bQXi+S6FspH1ehVDaXtduY40fi2PiDF4aoWkqNr/X6WWyeBwBJmhdv71ryd0sy4pU17gT8r3
wBxQ9GAUv6wWevBwqmZR/ZQpZQn98pxgBmmNNLpzIjQ/NoZa/LQk6rmnwIXHMImgVZnyCk/2GJYD
K7304bSRjcf0z1sIlOvD1GFfg+HifQwoJe1NwwKFdzVM0Bb4nLfv6GcL+R+0dQk9tDrx7/UgHBh+
Y0A4IUQbdL4nH4KKCcDuZ3558Cn66vx8GBP1DN9jshmhspJuZ7hT8/iN3REGXM3whJl/UnMCsyQO
58Z5gCLTFZVErmLLJeZAOSD4im9wz+O25ComoCCQCim3MG3DRW4prBzkMGSCTDsVVn56+C25h3C6
81WSfhUt+oXbaDRE1I4xAiKs5NTdGcTchNWTE0e+e03Bp4y8tJQTwEpX52jM33oCLpu8ZG0RiQA+
QvahDme0Flhniq0ul2YdFNVxfE3mf7hcKusbwrXI+z9OD5Bb4fa2JvfwHkvThzW0MWsestfOGJRq
7mEd7Bu4kPWtU1U3yLD5RCgJpkMgD0ooSGwHy4rlOumKGCLbZj6oroO1vtbHEX+Y5AssDAsBXLkk
U2XqisoWcVgGJbZa83SfsRM7kMCQS3bGXvqg21UQY2xSn7Prxwhqn/IMGUY2cUbzgHHrO1PdAJ1L
J/OjsGoeS2e/XfF89RA9wUvRiVJ7pTQDreT1lDJd45BRKnDf/Kp8V5nifRXyIfESJ79ummqN7Xrh
l4U4mTqdatCyTzT2m7Sq+E1iQjVYbO+VxOY3eJHCJXZ9Xl+6rI/30IPH7R+Hh4DSPp8Gn22sN4Xp
IEuG4zp6c7WeGlZMyuI+1RZtbPVpHZzRGPEVy2dIqxzDChs6+tmPEkoX/yNjntBA26rX23A6faQe
w4QP+sQ3+AJ7CEZVvh7n5qPqKHEnSxv+iCNav4pqEduumJvxeNlzLJWemQWLb1wclpnTWIpF2zop
uJfdxvXkR6Z88kxXAPGSGoVzj/CInY1WFv5OChAgeycWsJG2DdFw/QN7JuDNT3rwhBwFZe6GsV1R
3r9lrSsfbF0zF9Mrl4W2kDJMAFWyHnvWbXH2v7rBZ6cqfe7YJsF6hdtFEzDzsy7IH2uyiPoU+dUA
I/0YPmCcrDO3qLXcYwU1IK2154oo1gfoJ9lk6fkE7ZZm+CYlejcWujWDRk+ODuPuwohOLLgq1fzd
x15NQs6ujjYhunEt+V7/Y4N+k3MP6fY8RXfG/kfDf53OLZvRLdRXslfs8Nl1Z8aa0Zmyu5VhZrdL
/mHFQd6kMWFIOY6QNZMNExGQZyR5B0q+bxR2XATATgHpgKmVdkwUpfOr5U3USCYag4vtmkE19Zla
2YZBNp/PqTRjNn3U0tjTcHwxAMcbXxGqedyF0EKfUoFCI9Ac4MqoZ0nMc/aoehOgVmiUk8M+DAVr
py7LDHAT1p2iTJDKQqRGcarvpXb9YDi9aXLHisHqkTzQe3hAsJT7oMzCS3BIXSvwvRpYdHwYTJhr
WmYMvNxYhNpP4tzPamr35sc0IxclpH+2AGt0FeQbPj0GwxeUq1TRGHt4mLYZX1xKCO18607Rl9go
27JnzEs0M+qeJn7cDI4OTclomBcSQM+Fn0n946KwnjPdi30swiQqru/hQnB654JMLxsfDpNY9Obl
MunayViHgORPBnseTYRiG4e7eMS1LCnDcVWJtiLWrfwFK2KIts8wkx0fAXUvPNpi0xD4wKdxQlD2
OkeoiGLe8GE1B8J4gGo+itgnrkqoz+wZ6ZgRUZezsajZMs+aVAFCKPWt58g0ucx0Ssi/nbYlaPI5
6L6cHH2GgXMkyIj1rZE+oi5QXgiuDvRiHbKTWZsKDLFd+U1TW6SePy6D6FpTZvT3YexfRd/qMjAs
Hrv7qOHMHWQn+2N28MbPHDZmybxgyoUcD0TGPalFvcZ8M1gVsCA3qLLkDFVfdso/g7PG9OIk6rVu
stscjP34x3M7ztuBX2BXHhQipEpUfjg4DKuGp0P32RSaou5EE9sMICmt21+H2LJs/a8yZcZ4bYSr
MxGjEgEuUZO7RaFu9gzwC+jZc4h4jZ8WVvfJHUYBcPvo535pSPr1o9V5EI2LWg4wnyIqeZBJmZH0
0aBR8LOnNWD436zGPD2h4Ew3vuJ5Si+Rt/DbK3LPfeUMdJXo+6uasnFFuhFtSH3ZtcmvA8es+7mQ
r9KO8n/mPbrBrU+m7ltZDPFbYVvnvBSC/5dvMrSpq7Hu/Gj5MGyaAE123lGDCYuO4RKqRvaEhtWA
cC0AL9e3Tg1Eym3t8JYojyYOQ/SWqZWDtp75rVbdAw+ApbldRueXUYixEND0L4OeYr5sWIq0Tbs4
IFnsYcA8pdrN+ZMgOEceJ1ZBVycbID/mCMq6rp5De2AAMHiqmrZprwrguXwRrwPmC6AdjAq+C/Ln
aE0RWO18PyqkiSIc13X4PLD9CFXxcEEqZbike2GbU20dG9CPN2KuD/YfZaIYa023ZjWJRsaDe4UD
UjHNkSEAIqUxs0kKNeghvPc+SpMBHR52TsFtDwce2KbZBzl+itLRAAtXy9Q4JMfPRS/Yfq20tOg8
v6QWzlC7DyjkEBac2rvPf9EQZqJYgE7FAqvnLHBvwik+Fa29tL3upilj67J/bmGh7yf7GIKzj6YR
Jg1Y1wGqoK5ETGnl4p9KhNiVfGMVIDWIa9xrW7wCQtdUkxPA2Oizzllqr/5EcMdTsHULSlu8GOBx
Jmq0jnb6O8Xy3LQmgFVB9woxHs1ZpaOVCcr9Ch18i3iTsGFhHdOvmEEehD0HZbT+nDJuevZG0P+a
hPmGKU/ly1fqDF2XkHnbF99FztM+pdBVSTeKtBVH2eRy1zlbqLA/hRic9s0B1E0jbQDDmrOn37jy
CpbOdUHhD81cMz5mPkTpP5LPCGm6snfvRcSmbyr/SIRyCxDaXPb4VX+tzNTGTtjlEJ/RrJgOajDO
ZonEdmJC0WSKU4fb6UDPBFVxwK4cCdyuKBmiMxbtEN1YysX5URzBxgZQzrI6NCInNFo0kLrrO6lx
bAfgFMZt0C1D6/rcoquQ5+Xvdp+klcPRMISsHbxSkGRanhaxVojjXr/wWBEATBPbny8KW6v0W959
WJdkTD85N1FlDEDuWSfI87bCsMIelOmP5x/hCZ+7jOJWBUnUw452ceLK2QdrXLwc+9uw5d2DfZOA
IbCSYwIR78UQhISqsJhRDQmiUPaEbnkelN33qCsUjnCykpSKeXiJDj8FRWRA0jIMdUAcaud8VBwv
GZ9Dnj9TBocV4+syIyERbocLGFu/+yANW7TaxZ8m8UruC9YdyKXmM786weB+zUreeLT/QglhUVjn
SkQ9IEg7SChk+uRuu/XXgsx/+XDqEmj0B1MMge3LhGYhBUDN3tip8rmQ98CcDFmq6eZ5BwNWHCzs
gRG2ocKn0kxA4+EHN9fjTEMo2WqCEqlBGelstSfu3EvwqvHb9HGbdVR4Je1fWozi5u7m63+Vz0Jq
rkGnfwkPluvdJPGkrCwc1dx/1oMpQe0jxDzgbQPeLKhP06xoNBbc10owsZPKxWMgff06GaQo7tdx
OD/Fq4ufbFNhU8dv2PHxPuA6fS8cmXKtkEW6mVnx/enDM9vkZezQNvbJbdfpQto7UoIvqk0pbclW
zAg4wmbYGpkK1xxVrOHKui65rF0JPpdpRbItZQ+xfYSEVYBvLGzTMDnuXXG2G9LswUagkCxEjm35
08UebBMiSFMaJga3wrnHLGgRIRXaJSdeED8j1tjkoNJ3zhKUdRH/Ma+Mw+DsozvbodlPr+tVSFEF
zhyvlWV4jtBXXi+LSfoJZZCKPH31/qmtaxpzTUnlCSsoaYbldaWTjKPZJSXHyvSExo0Ensa9448t
FsGwE7VmmbxXX4O6n+wmz4axcb1ZF+64kxfJ6bTSgzNSoGddHHAhd24WVbg9wblv8YtMe8nvn7tP
u2v/H7seFZmrlGfTzf+CFnl8kaJe9lTSMu70RQ+++q53jOJJ06bpuuLuirSoSuZF3on7i4pxjCpX
Tr8L2wJXTTjH6z+hZ2uDkYnCtNAtgn7U++lnkygm2/BW3jC6vKlop5nZYF598MU2lrwIXzOedMuc
7xiwGmBJcyJVs7EIWABJv5WdBiZX4y5ui7GnOVJ6oRcOvRc13sbeppkY2fs1XYW05L+XHbZq2l4M
+ztdbP9qCdYRzJaWKuUc29kZMgkcbpUJ7VE5Q5Y4WEsKZW2LJgOOhPL8J0Dx8lA5gcHKZaF4OxYx
5U66FcoJV1pAvHVKYFUzGzpYqmeyftVaKl6vlQ1x1+RDa0B8PSSIMikgikhhSO76yTPLtVO9Y4FQ
Hies2Bc3NTXJcXoLgCkmNb5mhlj5bgL7WFmjv1kXry0Bxbq1NJ1l5S/RBfqq8TWIPhx0h7Vrzmf9
74Q0vinOfRbro6+u3QMa9w76GEwuz3zbkAiO2+uWr/QP51duL6kpDr5IIStEBG9vPFXvTnCJ0ASU
iNLflPMD2vTx7/2OWgVRUhJVcpAxgKDgKeSQnOH+7JafJsQ3/me0OS39D/1qVvHM2uEM6LFlrwYP
tgDFODFdy6m+sAS4h7dLOpTBZF2fQkER+HBaK5Sb+uWeT2mlOizWG3vRrFJW1q15UsHjHmDHZXTm
vpvXx5vFbhJC9QREAWoX+mZbs8kcK0i2n5n2N+42xs2SzKIVOJ2L26LhfWQ1K6YgfFmsnuwLULQ/
QuiVZXQ58Bu4TIffk5DnH+5L2GX7X7DsITqxI52MiR5ls6dajiCBOoiNu+h5VulOMiDLC0LPeano
1/4pioBZxaX+2RsUmdM/Cenl55BMNywpDPei39ZauPVCNehbeibzGyBFDpBnd5bNNL2fx0AUhwiI
gGojEMTXTfYST7lLc9q3ukoueq1YfvZSGx3zGKdz7eoA9uX1mgqZz1qL0xh28KgrzqH0jva/XYGf
cV+RhlW+L4Mqofd7PtGsDLOdfm4Q+FTawiFsnF82MUs/pU2r1RmPdXCyXIPBX5JucTaeUoB/4APr
ZaWPS9nNr3sOYrfi6pAzR/Farae02fG1FU+LlphA66u+Xh16WmveEUiVevXv6WceSz+Kj8uf79t9
QthlNhAhZsqfG6Pt2r2tPtkUIo+i7R6DsLx9Eqy/eK5LH7iSSvbOp1GYTIea6/WuBmGs7ikpPf8G
G2fzSJG42sQtEMI/SLgl9EXeWv1QriU+U2GM1Mlyzi5uhnyEAcFVpJ2Fy++lWmsMbT0OQY41i0PR
gRDMmINwGggBbkRfEcRRGEU+8RjgmlZBB2gdZ4XmOs9mO+FEUyS2t5zYplAv5gdAlYRAMzC6KYyV
msDh9V5QLf6c5R1rFx1RXi+MAZQF24Ed5ByqGYIeb662avRgDls7+Z8q0VlOOgEaiYPwBE2TDkLr
KV0KNf8VwKq2NuieV+7ii5OPJz78TaufYhRsnTWmSo4tRrmcNKoBZYysOkA/aNba3En8KmABfxOc
j7GdrvfqFWvSXRkSZ6LmD8ou8miaOyp0h4pn71sqt/4UzBzOoz/TA89UDugzk6aaVkj2XaLcl9YM
8Y3zk1aKq+udF9p4Gm2l9z1lOrG0w4wJqbid/pB54Vno8yRsbBdaeMCyLVCopwr7DNV3MHPSI+/X
liHhlr3O0/wvLSOkghQEnmjMD7zP8uISZd+3Db4j0+uxzWRnnRVH6yXGG6rpdt4CE9LD3EGFxv2L
cEbBOoFS+f90HTPNl3UxBxtgn0aqoy5FbJBGIGJCMQyTZMIyHKf6fSqpmf/SfxWTckwbhv9jIInE
4NeBkxVSV/eN6hIyRCDgsZGSqxc6hGpTfTO7l2xpgcqO6qC+lHayI6F5ngtnGyd/RlTTrf2uzckf
6Qd4+2FSpC79uSbiAuMivK11o9+G28c5NIt22EiB3EYsBd63KLvcgxu01caY28UC81auuA7dApAY
6mN7UZRXEECxVZ+FvgkPoCs9zdKeSZGCY7EercO6qw9Y3/cmUpWDNF52T+dTWiLXRQqBQVVb3yGh
VMvgEm8RfFeBvdbGg70PTsaKNhg0TZ2Lc2uMYEqflL42ku/D26Y7M/dlS3KQbiF1FT+gWgXKUVmY
6DDJD6voSubnvA1XAKYFJDjc7St/F7pXtFnDhD5VKvxMalWnohhRWDie7kz2bVaAjyeK88d3ZX5a
sx0F7VBHCYebMev/cRmOzehOsA9GWd43D/WbWj3JZJ3YSbQehRAVyNErhwCjoIBsEkQr+fgAxopa
GxTa6lRtjoLI+HW2YljhRuuOQhljVy/wAJyNk8+k31VNVrTd2quofrb6QL6sK+bJiyVojaY0CapM
ABgUT7OI7RdDzpTFD8fFhvpuRRaxCcVQ6QfECiBNViU0KO0Pq1R81VbK/9z6jmcaEMg9qH6dK2g1
eZDOV/kY6GDzCT2Z3VHEjVIKFGEc7xyk+LVFRMx9M+f9UVg19OlXUigbEE9hDIW2vcKov98QHrhy
p9awnQ+A7u/6inJkPDRROgSwxsvYdgQrfoFKnYGgMTKJpNM2THfeZZ5xYTC2DqrTFovMyllX6j5R
EUlXJcIgsd5Yf272Bslc3xRkotdIn3+7wUTrHgACjsntOLXJBSOBMz242PbzeuOoZ98DR90ZpHAZ
ifybJ7E8k1ylrr9BLN6FlsoODClEqKTYV7BA3JTBJ2nd2fcJah4y56zXdgBX0zOkamNQJZ1fDSHl
drKvoQXwp7N9VTip9LaLC0b2ffSZbZEn+fiqouzp5b0gNjMjAmHvQ/VPfxNQqJRM25KezIq2NVQR
1f3xaFA1iNC+IfpJXMMS2LHWXfphCm2dudEno5RXQ4tCV+H2tb31z5pt3njMnswqU9Geih7v7q1X
0BhWc1Z3JSeEQ9rdrcwcdweCGvR3oPgvuq8jHDWEBFmSC+Zg6kjZ4M5VR9ocb2PwsrTVzf+y6U9r
xo26MfwvGYcxS+62j60hAUJt1d/WvkTQhvLGH1L+8g5pvvGz3Hmj2LDnTRriY7aWXc5ZlKRAiw8k
0hg9W4ee7c2ApgdU61i6WAZ+QLPPx9Lot5sxm8ao6DdTaPgIdxMQLA7NEtz1bJBNLgsJkVxVfu+c
T0J+HVj0vR6J+J9l91xoOutsIjE+dZTLfhc7lyZKQAhTR2LLzGf06fUm2wOAfQY86wuT9EShsxrd
OfIKkOdYL7OMYfKSDXjOu4Zd4f3q9PwD+CdQH1DOakKPUrnpSe54OunZPGz79yVbHk1ZqySjkSzY
UToQ0auErdmIHHf2MHUKxfzeL4Qe7jasXuca42fakaI/SzZkA4VMaPGmPV6u02QubwMocqZhd0p5
LJaiJtioH03vBN3FXA3SdRQp8iBeHsUQ4uQHhurOB7SU9ck2L0rMfZ0LrqA3cVYcBKQHtFM+FYOl
9jW7G2/mHY7+eRtLBusr7wCpJyTCpabEo4gKfYYCaJTbPif6LkDrEiL5oSdLEPjL0KC2sQEvJGgV
mwumDuNa5v7n2BR+jV2CUMGII+EopQuhhu1oY+2nzmjAT9AT+KFdgKJy/yXK3wIBKk4iTCaBq73I
P4ia2qcOR046uHJH6gIbxu6kfVyT+AL6w9hCoG32gtiTaOrmRqMNFPQnWYollWEaM/J3d7H3pcmr
DQp9cFeazHXrqJSlFB07WegeP1wQ18HMIjpzBUAiMIcdDL1pYbFTLJbDYyagbC+RTgz7lsh1TXe8
Hi79eWRB6VlPKyy+nfY0UiOpwLE7scZuYgbNS085kbAjhyccWTx8e7U4qnVEbNvUqLAvIzCrLUMs
PRGYcKNJw1ok/S+XBh8Prygb8PVpPul8syD1HEFJexUfKeweRem8tlPn/NfbKRNmHfW4fP6s4Zit
VOD2nvmvWvSREA/Gm/o9S6YQ/pJ7c6rxrggvltl/UubrPGiPsRYek1ovPpgCbtLspyumSSb7vV+7
AhuKUy602DV7le60tZ8GAtanbMGql1XrkwAZwessObgKhLhXO96oBk0p5xBh30Lam5m1lQkJGVCa
v9ftJbeHDKd0DRRWi+6wakq8DD9/vgTKjnbhHriv2QVWn+gcun9pC7CIPIivAfTdUFvzkdnHs5H5
T+iSpn/Lx1jQ4eeYwocqvasKHYvtxRfVzLmS2JoQGIPTKxUCpA+XEmaVqpA9Ywr0DSF6MDrhvuQ/
9+s+5D7nI2v2y9jBag2itM6aMEKq9zzqwx2P7qd5PxJokPHnB0Gla6lZQfV0iJmr1dqEa6PONp/g
2si2g82Hg8XV0uRbqHw4uRMLz1wyfPiLcqOti6V+5qVhYW+08NJBOz0rutUK6XTFYIgjaE9Lb4Bo
H63M1VRYCa1Jm/CoXyeYIcm3c6ridNuOyitVqmF751+ovVfIjmHpS5j+pWQGMxm11oxspuaXkRD+
nQoZ6/QPIrClwlL3QGjOHm8DSU0p8jUZE4ZlP4j+4iBotypcrlWM7SD10anvun1Pj9dn1sNxtDF1
g5NBYvsCRQRXnQrWAYbSm88QDmRpilIFpBDkRU2G0nljxrNiYAZDSjjnuG9TPRdewCHY3LQo4vES
G/uVOFF78jT8ZXtQzfuR8ZrdNm5oRJ+TPMaRIOqIxs5YfFQav7mvPEEPT4IMROyEiRGPKEGZoRM3
+XkgHQpvQssBSa+z+YN87EcNQIky3LWMs7scM/ewB5XXeQEFhy4Yk+qWSCEzszHGdV5j+RKooXx3
U5+C/QeCg/c5NphZjUL/dXBlZwzyjK/0i8RY+UAxB6n8b1UZEIES4Tc8Nfc6tOWAAl2RuKDeUbnJ
DLsXfbipYY4OU0sh9nYEM1q/dME6WTY918HG6VC8pIwZ26yZnFvcKR2ACyYSTqW9Ylv3AUEQdzEo
QaKjypP811htKKcVF6aaNR8r/lzaGmF7yxHE7Vcfcc/b3UxAV+4f4lW7Nc17FWMbAoFUXCDNKmFc
66j4oV3dqAHewA+jYQDCjgyJuNc4ZkMv9rar+QvghPGdMrnph7hGDmTiQfR/RHVVDZC4OTHyAIBE
6S/4MzeKKpQGAy3s9ffxSIaCKWc8Z6/VIhBqHq7OVUnx5LL9eV0In+Lwhz++Lh6ciyYcm0o6F03U
lj/umLEr/kOkR3FFZl/48kJdYh2NDm/S4WzOzGyz+5VtDIBKIMsq6NA3nZ/4Vob/aHFV2ZdIsTbN
t17ZRaVx6vzT6Rqa/1672xWWONxnl2K/lRuHh5cslhgCBE7pfPrEoeg0RJLLjbP/7R1gZtspVZl8
23b+SaK6R46pZlDEq9U6WcqbCpNzkfXQHa4/465go/Ym89MmMyzwuFBNe/pKiSIRKJRR3uzC5SXK
/F2FGlGiIzRlZy1ptzGwGkl4LlnbTIIByjeumKf24nEtuxS95klxWOGeMB/ok37qGZ6hSlgDG8AZ
x4S++Ezp++eRLbuZlz5uWno1yX2ck2CEulo9vchSffj/KdSmkI4S4w9wPrx4cIDk7FsaL9ubZEex
8u1hMM6+kJrWjEFRInLN6aiLnjNduZRu+cOch++urA2MwtsnXqWEGv1asWkWppaTgY16b9lBr3xU
s+9cFhrmi46WiOce3KI/GxCey5+AowySB8jSo8HwdUcRyOr2DR5Og/rTD5RhfFYpOArbenLw9U29
2zp9lWj81l2vk54zx/wOTF5uMG0Juqmrd33DlUebdQ2RbZtUy8eg2UXwgrSDtqiywpe5+exw0EJ/
56/cXd7e/DdYScqhIxKjAdhb9y0Oql/DbggqyQxy+8Z1AD6u7LkJIrpdWjiavR/Om3IYaPrrI1N5
8+jUUWK/Aj1KWBxAKBa9m7phdwdeowmjEHvcAShMVqNbmckaqx9ObBYiPNQOdtYWeiGKGeJl/hhT
/L2b1uafhbOSSbJ44LInRUGj0iKMC9f8+yHYWdxTsiW7xRUvENKajR8jADh6LqQWDc2zSw1SyVEW
5tuSBmDmDFPQTH9c8FZ2VWtjWXnlbscTO3hSLWvapyKxY0YV/eztSh6o6Noy6P46I2RUajiONfBy
IhMGdFQaR9EAP2u5jh0XJSpdC76EUYeZlVzuwCicWhc69l9DtxU0DqbyRlsvndI71sZTVWpR26SH
0bhvgeUTrleAIWqIhqEuU49eIVRWoBuMbL2OHs5v21kLIJWglt8Xp7GZ/HMBbRFeLg5lMuTSZgUw
X5KYbCyM6y+hy5s8nrZMd7thuk88E8LzT10Q6tFY9kM8wqCHBXidl/CpaCsJ/PLSq6E8nw1MzgT2
RibjKQhb2dFCZQLc8/6RhAteyaoePimFwUuekBDhKRvEMtwBxaxflElksq+Y5rlP0BJmEcKE8S0d
k33mzhBvt9KNWB8C5qaqwuntBUVKEBcuRKi980LnLzZ7VHUOrGQn0qLnA0LBdXw0OFt+pyU1GVnB
Ka7fSASN+FC+LrxOsTz5W88nCPom82F+gORCkpI0W+JVYlwh95ANeZV2QT3zSTmfSVLTlqkNe7Vv
aUrf4olZXI0WiinCtCek4ek3h6iuB/wXKnLsp6xxnjr8QaHw/38y5nH3T/pbQ805h8mR5N3WvJLm
EUZU+ilSHPOfps1tnPC1JxxwdXVlxuI+Gjqpa38l6tfSmQ3JscguA7HWKsQIsqUeVWtgJzen0uzX
LMjzXCQ2N1ZO8X+uCeb/XP76F8DCcKwSbjkho+R6HIUdNtV5k8zPbp+Pkai/nNf+2VAYJCok1plW
q7bG7JsP6bAlWyhCYimrrHM/X9XwXGU8sAuEBIgDgyL7Xgpyk+mks0A0OrG1SiPfxwKTanC1sEYk
GOsqlwde5GZSc5UbGVtAan9VLri+k8HkYqA4e9Wy4niqUHCX3jRuQkOEfZEYAX/U4wSXBgnlywx2
pN6ltppb/Q708VewcAscBdFp9cwDk/7dR5gvAzKRL7ftIlobhLKsq3Y1LkEgkc4Jl3lfvGZlZevq
dIyy59G2hLngO8YtJDfu1qtwW16qy5F3eAZnBZBEQEhN/DMOSucUbEfO6CvQ/k2xFYP2g/YxM5zd
YzPT3jOcyuZdjd206Apt03bYyoFuovMIBcqpKs1gcw+3QpGAtSEtyaf6FyEsQHFgVP6F79A1Mszs
obg9PnhO7Vx4+xUaq0T3A0dH9yXYKiFroAEvYJPaDXbpb3BMRjG5z8nfiO+qU4pphmk79K3vSaoM
j3NBjLMbBX2l/ZGT/KI9cUpZl8aix6fEqrJVoBrRTnXaLSRedIGjTJytv1QklBheNAHpKi4kK9ZZ
np7pxdKrLwucJohri5GXn3PWWezqiz3WkT24VqYjNsNpncM+NyLBcvLaUcqLx6ZReNt9TWTZlq50
MM7UlLUcjhDB9jHgi6n3GmGd5+tLGv7dGE8HTSXjTTwqJBOdoMlW98hlzWcQvB6nOmJnWDbMIf4m
uqJHvEdCbpmKYUT/8OFGPi2FoNFAGIuuYs0iRAtwTJrPRf3B5/2aTEY8FcaD85GhdEjwG1HkDO/1
BBSBWDEI88utIqbD7g4cpigHdnGDAcWvMP9A4gQL0end4+5DHx7ekYsV32rCQZfBmXF+j/89/QaZ
HKmHhEQz1GNUE/JQbb8Dq+N1cRH1kpzuiIdFhOw6zI/AQ0Ix78OkOdtJnC5Ep4bWFkKuJkiEJOxZ
Px1poUa9MYJr48eFymSFrLTs0MadpRhLyY/kQEnKN7pM6NHyAJDCXUloReM4bVpKOU3zPyPbqsme
kThFwfMU9QW+4Y70mGTnFJA/6rIRMMaPBEXt3C+3Mbb1aQI6uP9G3m7hTtOJ/2IB7Za1RvGrf6+G
C57yo4FBGIAAgYcdicF4dVEUpn63QyjLHBS7DY8FjX9oebonFNZXzdJMq2xOjOpZSXinZngkPsss
djebCFNwTqFOZJ2Hxo+ZrVmZKFYOsYoFQdQexhw+E/tskzR9fmuoX+K5wzN3IF3aHiivpijkmJc7
yUiA0Uha7hQoLGyLkMq9kqLiz0G6x7W43jTAQMiNlDfhK0uS3HA7MZbUEEJbN3149U0NgpbeWLjd
MbNMsEYvoBoTruexwiRxX95lVUyxCgyLXvzl1ZRkSuWZqmjZY8djwmtXvR2EWOshQa+K5I5zU25l
MdRXRZWmYas6QaVSb4QmcHdraZU59mfoRFMuotspChkSkQDT5C6Fv2HXkWLB3a/mw9zg2ZokIhUF
IItNBNC0JPQILcw//oytbykHWOXA6tnNdLlBzH+QJwaQIIQAIkedWWy8l5PlFuPbChGjkXksihLd
NsMrVPISQgqlR7AaTUbM4m5UDJnA9TKZWbFzgBEUsvlHhQzkzMt6qqDn/VuyRjbXXodndaWB1Tf0
eni9bGvwxrDcQ3JzJrBm3DV4MALcn3TIR2M4amlhjcQv99pbkBuh5lFNsr3OoMVb101gdOqf3zg5
F1y2QMX/ayBHQ7LIF79gjRO6HR7eOgNh6FIyYjnr4sGyD9yTaBBNDRVVHxStVPOgikJIE3eQboHm
q12GTnt9t8t47ewMCthV2fvCc0wbDTnte84bvE4HcPaNVMdSkD7rgFZF29uiCIqbRh3g180nruX1
tyMQpa1Xl++SmS7QTlKALe7uOzKG8+QS13RtT6keOwbHj9Rcp1Jk272hcTRV+vIFJczXXseZolPw
HydB1ypi78HxoOD+NSAJqn80DNu1zEnfzQGrfEYzMkN7NjvTQp2+V39uvksy2x6auadYLLP7A5AG
vMwCH8NcU17MqMrlW3pu02OCMJfacmIMs7/jc0TUD6BmDQ8UOWKYXChD6Auoz1yL7roAeVOikOKq
EWQPbfa9uzO+29W7WB52PBX15G7dbl4jX93z/2LVWOavjadnOVDBX78GqiaafcJUWjgalP1QJOp3
bYeNcu5crzAxeadu+e1pmCWmwD/2c9pJkaNWlv/x5TFKp9ZgQVG0BzeUtCLj+Ysr7aUx2W4Ht6Zg
u3tjeMVbUS47WtGAfKTNc1797o6WGDZRrVscostFrdUnDTyM+aoJWmYND39wPnp1QReVJ3CCQvEf
IWVLjk0alH3ZAgxLzTohX1uKRSGfZkTaVFvwfNwWAZeVoH5CeQIC2QDZub+glprJYkMCC6DlEYPv
TVYBVtyEplvEeJ6bjXlTdn99PvTY8XKwcmE5MXZ4jmxoDbYWqdQ0wNDqa5EvFpDbN4PXVAjpY0Lj
h/aBQ0WwVmtbT6Bjcf91aGXbJUwrpx0PBqOeRWwAZwfu4XQj1d3m1utoVcJqtqtci4dfrFubueRg
dlO7wgjUfRwlVvUv9oC02enNwoXalFaZMMBlwTEfBEgpsmSC2i2FoOTBQC2OEs1kva29t9A6QBsp
Zw8d1ZfydSpkJdnbS8p5Ezffc5OhitiK9jtUhZuNSyNkU/lduEjTZfq+AorOebDtnqsNM/uRIXsg
X8W5YoR86aVEAWctGm5epZgQV1yNkyNbEO8hzS7TWSCbs/zPP/7vmo8wHt/g7Y/rFXvFiwyC1aIE
3G2OW5Kj7chB5z4C4GbTc1r4BawYn0VcSNIvo8ZwkeY09BTAh72oTtzi57fKt1YxsaSMLxtxwSm7
Soep3R6BKGx7AkKB9VNX+J+O6qbVW0MrBAq+eFmWZVPLQt7ImqSAa5jiAGcFgjK79r+vuNYVTXKj
xIsccMtrP1q8GjzFGL4W+QnQKwFYFzWDXiP3a8xO1fNhSFKbc1Lpm+4XhyLenLZ4lB49AjLne97g
goQn9inHOFpkroCWwHheGTRgf12YTLam1SNAf44XTpJLxYGvTutZj8MDTejsXbduBoBDz6Aeprd6
vmuslY/2OlAWrK4fTNqcv4Fq8qQOjrQI9lwOHD6bheTDs96lgeM5LKEYlilDHMBiVXfa/eQpzNRG
uH4TyQffO/kMfIy9FhhbaCtHM3zL+zFFgg1LFlUud+WibwFjc/T6MqGndFBUz4ibnjvKszZ561vG
xpu2toyWA6GWnYA9Kx3ONVfizJ/kEK6p3MU4S5ArYyaj+KMm3d+h2W1QdUCTehSaowXv3ptkiP3c
e6IZ8ib/Diy7AGXjmeSl49j1gTsa/GwWkTdVUWaFfen6hmI5sma8/91lUBvvotUNRFSZNU6zFufn
YZ4CuT9oU6VOnY/6R+3gKBmopDOPJkP6oPvlwqhJYQqu01d+J3koV9fNjiNaoqn0Zh4Znh6IRTiH
bTp7jz1EY1+bUN1UFDOxMF5msF/+b/mmou4TlHjbxDvPOMNlVFvm5mR39HlymRA25HRkg6KbFqHm
DEn5M3ApQahQn8NAo3/efvJ9SzPYnwdNTZdWi+3WF0V0yhi1q1NQEs6r1aAuh1dFeYY/5KAkWKQ/
QPQSOXow9gTtMt5FsGwhFGhMU91fw5WoM4pn9096gDBgXidZvm4PuP0GD1PylnI+yxEscIP6NV8V
y/MALL1leo4CbpT+vmqsB4VjKQo1+NbsqZngO4iJJZleYFwA2ihDxx7D5y/mgn97OZQX9j+D0T7d
vmntCBs5/5epCqE4sl1uU29YNAyUE8zDy5Xv5351DW+JgdHvcZ4AaYp7tL7S/mPISch1l9xY7sDc
yPE9IkKyTPd+B2KB4fqEpYZ1MoQv1ZJkL9uLZKyA5mq6brrWKVaC6KLm54XYUnq4C+C2+2k92D9P
YYkrmE/+J2C7k71GTBrcbkLsO7YRMeSxn58JyRJx6lbssmmgdpDlVGIOfCordjE9qvP9F7MZeWdB
XO9shJz8JTlCbCNc5J/xiKF9U1OOKkDqtIIuSnqE+2RDEgo8bzwbBXi/MHtMBrdtuQFALEJGCpvX
YpsEJnJJQc9bjAvE8DrSjwCB0YiLRn4FOR21Gg10gv9Dm1r5nsemz2OJ4LTIlMjP4mF110a3xAbe
A0F9Zk9F9z8C/l5emTaGHRNzo3r5IOVJiH9x+xlrj58OCdL6zy6jfXXXnlE0gJNihMJ0oSQ8YIcW
0u42hGLdOtT2XGSB8iB+AgppKVVroDX2ayplGFv6Vas+vtmyvsaVVMDLsHxLfHKYk95Xi0gHCFNn
HToqxW0Gw7fOVsChm5NJCCRcMJpRIbTydZiaXpwJ+E1QTmM+IoIQW0PSlQu26GbvvfwRvkHjlV5j
ExJOr3TPEd3ysQH2hcB5S61MdxC1tJ9bkXh7e5H7ZvxHxdEGLTIM5POatZ3ZUG9F5GrmUwzwBuKU
URSbrVtt4x2ADjHExhc3c9lnSVVd8gQV2Ju1UuJMdvJbhbfEHvr1BctiNKK2MbnckMdVtvBjUEpw
cacwW5L6kahe+S4vvJfmmjPOrVPTF0xR54TM2zXc/Na3Gy3hKvHdq1re5ClZC57NYKtiaiSAOIUp
B2ef7mUvkjtO6flnTqZROvYjPa0XzR3Yi7fyYkBjUzRp699ERkgiYCo2hGxuHJ5BJUT/A0Z4l+1+
YLMQa2TP9xwxZA/D8itviILoA/IwNAhTlLm1oUK3ZeuaJFUzNHfZ+aYDRSM0TZG0br1jMRBjHgoZ
FGhiKRT7kXEC/kdB67AwhgLu7zLLdTjF7kTriSL1HHENfB1ImVv5wMuRW+y998aO7mVQCQCsvIFM
+GYrZT4t+VwIUYHaHPbP0HIPU8AyCadZuxUY2rGt9OFZrmkvyPOc+ex+s0LG8j69mi3g3WI89xnT
4+gFJFNudtO8XXWQ+0cdzwYiMnwHTJ2FGtBM2c/NBTmaMZLXdNoGcln20Ufs8EZvd4CbmAgpxI8W
GzhMHufWvxXZMUOFDJvHYofLOiuc4uvjkb1MyLOq676zbC4NsehqQ/77tckUIWdBv3c+eNHSm5sr
fScSAi4lpwi2hjxRngSOCAo8F5WMGEv1mv/TfAtdDPIkxoRfWXnMekILU2FYxN0c3ECR4cuyIzaT
pUhiMW18mtZXkb7k2DgFsSbx1d2G6ymubQQpWwl71eg2jS28dCx9arucsK4k41MxKVSL6prF4UpQ
7/7ZB0SVyp1vkj7DsrjutANKsxqHDrci7RuI9FAVZUA/qz++/fPlk8w1MqAIvJFztgV4Mz/Ze379
zM1CEHYq36qQo+lMie+iORqql8oauuSVO8Y4fOfW26/0Pt0B+gV9r5vSDgA7aMD0nJxqtlSpH0Qm
Y5lfZIUW2aE7X0tBQ2BxiFR7pSZSd9karycqPPRujKakvtt3XQl/hkNFIVuzt9p/kKqikIUQDtbD
ttNcML1Yc6IDLJmwJ7snD/TC9dhLI5qqSbUcBEPdR/8bFV5aeN9r2Dg10yQgDZGNebwUO/UaXNpv
N45YB467Kgg94JEq2Wh/v6hDmRpmGXlkCpkSOmqHMCtGh/fFJsewrMqE9gYTHtpzztWjoqZ5ZIrj
5RW7Ho4xsyPDs7i1U/NhTIRpA1OmhNFR6i+myUCEgKvVnngSQCDl2qss+b0CWKgCO+aStjJ68DBn
xtxOJue5mF4ckMKWpK9sMYSV2sYaKdLNqU7UpcsbhO2B/6M5AU82w/yuSUTX85sRZ8SRiZOY+sa3
GT+IzaWGQUJ0HF6fE8D6Rk0B9ojMV5I9gdW/elFuZPApk8aw9B8AJyldPDU1IKSpOB9CCs+i+aHr
BA5uIaBMuWUNm+RrE4+/YwfXSwwWEkNFPmLnM/WXYFAYbkdqhGHv+pnaNIWSlH3ag+tHtnhaT2ac
b7FEbPFqiRPrdSe3T7pbeb/IwNlarIcXdRWo6paXekSWz8/UN7zVbGFBW3pEsVBCaaB2AtzfoP2T
Lwk/CJ07a4WaKq1t1HPNYfpkhB5PH3XP3KoSrwHlvDV0H+FUqACcpNIbtNH/zns2uPN0unWeyUIq
57Z391McpXmIhlaHzvlPI5aPVjjhqEM9M76gb+Hgw74GSZ4MHdtIKWdcWXl3g1SJpJn5hdSGS6lh
MS36kS7BsO2JYNplosJ5WgWYNTQgS4hWRA2/9VDbIv8+szW6dSBIttPgAbT11KlNQ3pp2VD/PBBw
h2BEAKhKUa9AMUjd4mbJ22/6fMydAeBEnUPFxrSIhaTewnZT+wNs3jnKuJoRrTzdNtb68JTcP1nP
o+Wt+Afkkr1iAbTZNsZgyLhr05E0vMj6OkESPk8OKwqO6vP9ZG6nhQsrpqF79S5qBAK66N4u3W+K
M0pg+0lSR/PBYq5gVuj6R7iQkVU/7ovZ8J0L7dnqPFSsmSTcJt5MKgin42GH8Udb9uLtO2QiUqLt
Ew+AstydIl6UbJSB+CfFdLwWVlZa8/ldYFViFoJXZdpbWxizz1vBCH8mjZRLeGzJN7MqpnEe8wF4
Tb3qt1rfgcFZgsV4MPbdsgeD54xIJH9dpMHSAuFry12ayWNOplvvyGYOsn0Tc+oV0skG9szCzJwj
3X1gztOk5YJNU/E23Ibqj4Oj6dkXpI90jJR94Ax5mGztBX6dqdHuQWAW1fnwDOVTXMAeJu0wFNkY
tkBvbp0e2ZQg4RUGfWhh24a7sYHS3WkxVUrn3Dw3KIQBQnUMFO/luRxQrOi4Qu90y1Nwyjtk45sQ
R/X2lzCprd5VVTYSaDLq72VM86gI3SALYM3cHT+VpobznKtUq+0Na1OpXA4pA81SSwG2+0AlFlhe
zROBlbmPcwFLTLjFA/eiNw5twYVVw7L5k8I4iUIGZwyWYv3VBASu6dY4BRkwHDGPhLDMmS/45CiQ
xpaJgGNBxnf7VHZE55XzD+Fgtmru+lwfp2/cyU2uB7r/qRbpUK6KQjr44WsEPn5W/84IlfGIpKTU
Ya8CBtjm1p57aU/yqZIUZuBMDXTEr0Ag/8DY3jkCU7ciVNmUImn68z6wqf+uLeCOu2eRS5v1gBn5
BCZioiLbLBXtfP4ImAKZthjUuIvKmqB1LrcZCSccFF2PckX0kOkD5yOtdw30NaIoJeKELsq4F6tU
cipZ72fHkl0mkCtLTS3FL3JSotzKLd6fIQwVq/r9xE9aaH59qTaKW81+gBcKHO8i1hN6SFbuKquQ
/iV380hOZIOTvghu5ksiTSwZZYoSJMM6pOqYc2IGXEnxjIBodLDc1YcM2ow3E/0aQMFsPA2JDOce
jlgvplTdj2zLI2BRdqz6V9w0/0OU7IDzF8MSiOa9vYQ3WMFVRzwyrNx/NajDx+hoSNjRj2n/FdnR
IWUsPeKwMrHpKvDfDmf01uXLf5KZGfGHXkRmvB8uE1AjNUXabPxcB/qJZsK9WbbUy2Q3saR2i+ZT
1V5XZDryVg7qqY9uDbaVkyiFPCLm6ugFOEwaqObda/auyhQdLDuahtQVSi4W+r2fld60qvsqBpKp
gKcrAWV8Qp+sSAZvaCryqNQNr6FB699cIykE3DfySGAKJ7S0l5SVIgtIzPjRHe3HpCPiWZ8JzSXr
o4NNkLm7fZUJpUabCmmB85496Vf/f2ONc8GjpFeYLnicwbTKf2fXUMQZmHx1wJesI048CQG3mF0m
mo80y04EfLUigM2oTdusTcFNqzetlWJz5PmR7lfxnpV5Pz5J+zP3jH4vTvvadi4OKbWKHfXdx3ho
B45kIRKLZj87h3jRpiqgR1iI8yZWPDlHhxBFkRPFu8bP8Fux3apsNgk/7r4KqTIJ2qqKW75cPOyE
OQ544DO/H/Y8ejY3ISd63VaL7Xx8AiC4mHSzfOD2w1r7jxS3s2i++BXqKQ+BTndDJL5MHXzuPogO
H8zycTXENGoeo4e3ZCQHQvT46kHYilbJOgczGBmkdCfaQCe7PNaZY5iMfDTFqEREVT8FGyD3yjf/
VLxR7FqbVuJXt27mPXASxZd95kNYk2osuC4cH0mhTCrt7wR9Lc4UhFsn6QdEdZC0TA/xGR5zGc3c
eoLOpRCPcSoCkf83iup2MP3/uQMrjhX2Iraxgltb/bXMuzKb4ZPV+140r88wjORstQlROZvMC2u+
cKfytDbkDJ/McunVpS4YZZdweau4Nw8hhUsSxj+6QGnxeriYt8hSC4xWF6iOj6U7PL/q0+Q4LQzF
jxFHb3u+SCiOiCGoOj/G0J27E1yigVAz9gvvp6aAob6SRyyYNIZ5V7UlpL+Jm07fQdkBpiZ1M45I
r9wZ6XLrwl+wuiGdo+PGiVpLGDL36VaQCOnn5e+78fyPKPmiSKusungD1rsrbxdjtVtvUtHl8Eeh
L90fckbXi9+88J4QKkBjSjJwg897hjeFLiCjzZjH+Coez1AtHrVIvbKserwzXpCzD/0Ak/G0IYmG
zBW7vHP0K5tPIPqVAoejmHAKPY4xu300WBLdEHmaGDvTHFmE0iqnwzrBGSUOsqjdpF5IRo9mx3A7
pIW6TrfltHI31g1rtbI2ByjUuEoDCoNOWaResWQWTGRurX3Wj8ZnuwW+n/N9aoLkZ1MbTGiD0wT/
DykEm26unbYvj3CWFfwvljfBpF+s2Hi0TFZ+UcOBweIIKhQ1jI5eIudASvJILRdQtREL2YzzCZTn
t+mZxCKiMYDsG+CAaY0VybO3SUvoxlQe8csvaqPYLS/04QBszdkJDKrESs3S3fMxC+XTupW+RpHG
AQw4m35U0d0Pan0CD907qEzPsLk6n3/Fvwa46lX81sT/kD3tMj/ba6F5hrW9ucAsp87sGLXyeEh5
oIbF15p6SmzJWbuYSUbqk2Kpx5XqrVvargf/rDXpjoHsmdTk99AenAUllV8MAl8IVmzSEL36ejfF
5JHX/2cPobGyehdXYeBpmja7LjHELCk9Y97k/2DTOjI++Ch6o1JScOg03VY5xUhqSHHCe10x/6Pn
hstK4+Uz5104fBpTo5IJGTJBXxf1Ir6M3ksNsY6YwrmKIubBLDV8OTy35YuhcAbi6CpEkUTC73GW
48ZWucZX5ujs/Ssz4ej5vyEUyHMkM7GF3vBOxzC+aOjdktXX5c9FIdhlXtrnCD6lN8r9WGCPHoBY
40n1cbUOvC6ZmRLtqnmzAHmFNuzO391N1MUiNY2LfO83W2zqkCxqJMjgvjX8BVnZA6Pdro4ujucc
XpljZh8M1CEF2EyYWZ2sx2n5jwBycffsreFSSYTpTQJbF4yAqZ3tBQfXie7ytQw913Qb8gy/lY4R
xQvP+Fg9bECP/m+2JFqNeq2UoQ5qEMsOognlvYiX8DWzXauyfp3wCIKJjiEWqp20p3ZOZkbEed0x
P1X4uBT1D9+1wecOqhTEmM/a3gmkyNIZUkPo7tzWSMhBEzAwIK2KZxqqzvRrL4/iFL87TLFLWWIk
IkKquha+U6TRnxZGUoPhsrimsQErW5ysDbAalTJ64dajK48tR2GtnhWC19U9FRI9pN3DVLRFYhcp
X9e9/Pm5p1XeaaaoVKXvkDhukmkYmpUI4RtUA6r4BiZdvf/rqibcjC6BJIX+xItVodJ9FdPe7kn4
iARjM9nTV8TAh6vRKQIVwA5vIopLvvv1tiU8lwf3bvAlcQR7Ts1+cYfpsysAhLkAEBqUdxXx+hcj
RNZDULKkL5tI7lTKsv9Qhb7LToI9nz4aOTBCHWxgP6G3Bi8gsKxz45n3iTBtbHLcJnigLMfF7WL6
xq+0YdMbWJBNRFBa4sO31X2q4+wX3iYgtr+RYZTMl4qLzGgmtv2g60dfBIx1uos612NLAgQkYv/Y
kWRmmqHL6PY0YdRe+wxuhJoLVu+mvzYO+Dgh3qM6X3eZeEkYdYtvscs3tn8/ydZvn9pMZ1E5oXCZ
8YuUFXyb47VvKGC+rtqkyfMtbN0oAU9O7cDffPyrhxyJJTng2lib5/6FuDy1CvYnPuZ9+8PkhuBi
gLoWApT+s0+TFX0Rq8MQ6WzMkItS16V73IALu20wziwnpm3e3BNwW1VfF9xrLcQJcrBxDt/ex7h1
eGQN/7ZnKDIy5rnrM2G0zplHpjeH3jVY4+cmd/yN60ZaYK+vFUije71D/IlclSH9c6a6ATUwbD9G
QuIykj8r9YG06Z/p+9I2zANZJ4Kg/m9Gd2yKq9W33Z5PWl7vgTU27ZT23oiL7MPILCfB9HyiRb2b
IosXQelkONB3WgY7B3gluvs/YHcKRSbGWM4rNChkDu2+1lvoo0GdNxGGEnGsZNm7lhSHwFKnSjcX
ioScm+MUoSxWF07oPn0mkpBa8OX/W8/CUWnAq2Pj4Uf4a1DhIIWtn2cMJNrDxwhSrEHPjCcT1GGV
5ri6EesnKjrQDD6kWJZyAmGM08O9Lw35OeWfiPDV1YUIyB2tvF0B6dkZU2DGhTE4mOiWlGZ8SKJt
SHuoY6cTWhlBwSwNcxeuUVxspT+kyXo1kPne2RBBYLzVBrTV/35tOWEJ41QZFBPMejmN9CvrgaHS
4h9hn28Gf+Y21QTYUIekbIe9seBkFJdVVLz0aqTYCIBu/dxwQsG+RabJGCz4prio0dNzdt7u4utk
8c+XN0KuJL6v2loRBwuqD4dNFNhBE3mv872z+HP6KUusY0Y8x5lAuJE6l//a5v9a9j8U0eb1W/Xc
ofQkhcKfjIoV2m4Umchk4BzDGfqZn5qctO1XI2MBJAkG1HIZpELj91i1/3GK85pkzZhYCVrPaAZn
1euy8r9zsIkREfW03ODpi5D9yNUBPm3ZmgNsii5WgMXKfYA+GK5+dHL10MJc5Dgz6N4y52oymSJR
nGukjY/XsQABMlHqOZbkIl5d0f+Vy6gH4ikPmRpvv4kqDvi34Ib9adXLcbmdj1RR+HSEPkZwSgBT
6ktPvh7GhFlqSCfNcY9HcX/xI07v1JWBBDlnhp96aBBVc4gkSl94/w7GsgQXhv+RZunI+RCr1y8K
CTX3a1WKyrheiMwFgZmlfQMnMT48H3WE/M1utAaO3mXlY/+ad0qtl+g1aLIpna9be9pJuFNg5sMa
p5FsamF7NAhga5F9jLYEDNeBgYOXv0PK8VMFKJwskeklHWawvLYbuZo2Utyw4v8dRHZ+/Y9JfYix
1zhsTJiSwSz3qyQg+JJhrWA9lssOxXez8oD5VbicuWk5gNJKXUhM2SNpoLz62Z6d+9x8PBn9L+6a
YFBiJ4C/pi2x628M3u60WGM+gOo7534IMwdMEekXg9Lkg3Dzg5KBEm+PZuQ8iHhsrCAHhL2t9G3u
q2bt9e4kv4A2FqB1g+B7B1rA4EFqGgHfQrJfBhdVuscF6cdxkKggMDEqFyWipiKhJ4+Yq21nS/Vk
xrDG3QXcgZYh/uPrTQzhDVZJVRTCE/CnMsJVBYv/WcrKcsh8hWRqbg3gdzKAI4RkhU57u+lNggCb
njtTQLoykt4QDlknn+ambRGPGED/nDqlaWhzJvb0Re1Rm5Trf/OF0XYeXAInbS1kEuC7oJu0b6KF
EUg/g7eLSjFq17kn7+HNptitw50tYHFPuOJbJoKIiJW9ug4f6Olkn17g8WBDcwNzgDaU8BObwjg/
YT5h5v5zLM2FmK527OZObNJjQHMRXA5iiWB7o7st+7kqVQ6mTYjRlA2JkTq39IgrsXW0htOeZBAJ
vnMlHwY9DhYaPg3S04958A1btE3MCANG7zdgJSapROqW5yAUmM9NTzSWBDQx/dhTKXKsZ0DhlAnJ
u3yb9zAQ9MndlLntZguGj8RVeXQaPtwxO+njXjbq3N5OSMEe62jJKbrnMwH0t0iLDeaTThPXDFue
OAOxkQ7k+kfD1qXCuK8GwccInz5mfsOxv1X+ycdDcJd1hNSLy46bJCZJkdpQoJUo/ofGlT4o+3nN
Pms7T1drRu0zLMrfwKD0uD8S2KeghwVbGwxfaO7k+xtkrulwcedB8BPKVFE00105wS6ksbEPD+pc
5BRLmkAHHhqdy37/0QV7XudOlU8j+RrE0VCtNflqVR+5p34HtpLHd+Tx9FWV99DqJJjPLCbLDxhw
4e8DCdUjruYm27zD/9+LOEX+8x8ML4n/LlXYWPVOOf/8Zl2vX3xFQckSTRNoPvFCpxvOknobPhhL
6xAyge1lbrIqqhQRjGfSzmzKWb3PwZLilusHvo1LI07UapWwWqK2tPWaigZCV3RrCK72vB7/yeLO
JebBPwQk6WsAp0jbF4/bJ3IUxhkrjyrLLf6zpUfbj179KgkPpvzfrylttyuHI8Dw/OAbqvRM+bmK
UAVh3LvebMCnpnNeDk4KDwBD284wIU0snYi1B8uW8Npk2Mj0KQph7vh77gDkYRNVwFzIbP8l3yTs
McdQ/aMbNmRP5SRKH7SlrcTOFddIz6buT6r7wBOSjqR7dCy+BkU+cDm/s4V8phijvQP7FOLNzwpB
TfVeTK1onXDlYKvKWS1Uls0A0jXiZDuSI1tuEXQq7kKyndBSdydyLmNTv/ylj7uFaJ1eVERE+41g
2YTStNeEnQiIp/5mpTmDBReTn08Q+RwmB+WAWofjuYL5J19EWRX+u0DIORhWSjNTmJEk1ewdYouK
iJaS5eVWN9N1wIyRpjNDR/+6E0D3EKpsC4haQ+Bu1/xc/PAyhp64lA7uoaIuUFsQnpnCW3qxO2Oz
FTZjizvD/cNIDDlMrMAPv16vkA4hVhyi5DzZf7z9osfJiRhPF3Kb+0TvrFSGIKffWqqfTrhLWHdg
p0gn0mux9gF+vsqA9KOciZIwRmytXV0n/7aerrwuk3H0g5Kw0aPSaF2tVq0O3W9/r8eK1kkLBVaa
kgxwrC4672Na7sRyak1fu/+3H0nW+VazTJ3rlzVCzVqbzpzP+URM+Imki4jEpzrP7zclnqMbcuKP
uqGI976Ea9htUV7WLVYOcsiL6GtnBMZTDvZ28xLZy9jfe4JGmCyGAJkxyZHZ+T7a8TxUCHwkt5AJ
u+7eTojuxoVHFstQ9y1a0NbZEtmfKPhJO+cgGkoexR55kqAOg6TV4MMWkPACSs13UIjycg0wzLjA
E2Gc7upiEAQNrc8dL04eKy1JYgS/HKmJD7yabmE+JqksnSHM19c/ELC6S+kHJTkMzOy8CZR1HIcq
jiuu//WN+JXfxNxAF/k4RFtF55sVy6d6AvoYVh3u+DDq8oL9/o9CQCBlI0JL0ho6rTDF9Gji4uDs
sj7wvgKy/mnUIYt4isSLzcCOwMBmc3mv9orrz0INZjTNbXQI3WNEvR8++6/0gaPQpPcKWmeZ1aGM
JLb09X1VM3HGtkTSkBzP1plSJ1c1Izun2XpDwcFPLmjs/bosE6yadcaVm+4FWMSqix7/mHST8ouR
chWQytvIOy1nRmHkHuR9kqffhzqhe5NbtwLSdoLdyozazwzHamCGtO9IFDIG5/Q1UnI27Wc9CihV
uQ5VPyMbhDnMcNpanq+lQNZH+iuUzWcG+AH1VZG/u7bddVEC/GLgukqO35y8o8wM23jPyI1PcmJh
MhsZIvARSjF+F01gE+jzDM9QKRu7ICFmgTqtmHBgIOPtSNXP+IVWjzhpdwpJDOYsKrpCk4OChJLr
wEVHA/M+9by0OyBqB7mgvq/lDRiC3A1IYeMvHgMyCIAuXSfB9h5H97RSy2B+IJSVKnatIAUVsjGp
Ve0cLMfb7qXkr8MoD1n3pssG868VtE3shvSMr0d0tjvIvc+k5XUCe9tHrOS9GB16HUeBQHtzzhU+
wpfvhK4Pnjoxux30jwaSFOamwqQLKDTrOcdALlZ3QkQKvpfxuuvVrBVg0zKMBhM2vKR9WcVMI1xz
TVMy6XyNrNNuTrF2Tg2/KwbQNDHaI0L0jzmeVUTRJiL8eRva7TSzbn3QGLqiMK5zI8jclXTw+BqX
3YgjjwgWSsH29OgOabZ52/UqDRnrq7hWb22hTT634XxdlhiODz4+I1tk78FtFyBWgMi839mVxYUb
/ZRovhYva+UWQ3P4UZ6hm8ba7yQeU8S7CCfPFAwBsjcMwF4SK125hKxr0p6rD9jdGH7KEEo7FNnf
1ywBLy604yYILjPrsC/gXov5ij+JprZj/+I/UvqwpTgikgURpY/uVVV5wtpef45ju2CBz7Gmzw6Q
n4M2BgbFYmi6r6Dbwl7OYW96lAelMYrHiJpEfpI5mOvsp8CKPJfaHPgeFK8VhbMNmNc5wEXBlETq
EuaOkgG3giZzdBWA2vw7RGiF4dhWeymNBxP/Gw0y03d46IGc4oGQJfn38taIHSAtW+HHPczuhrxx
eA3caC+S51fHd5UoB7ZkMXgZyGiF8Y1CHCt/kwOlYSsHNPfKsQcU52o9D8aAOLAqAhAem1eJcXH9
8iVTm8fWK63CRU0GCKM6j6fK+pxOSTtYRq6Ro1JmcqpzN6wfryvcPDZ61AC3G0o7yq8wIKt1t6f6
Q2xRb2UV5IMCKGyMfdUskXfriOggIADE9XsQszsKlCVEargJV7nU0YJhR5r2TU5WfKeIi9ciLv7+
kVgk5eyOtjzjptcKmBtXfQyCr2wKB74tRkKNtD7UXIxTHwzcs2F5cX8YkqTeDatripAfOxbn3QC+
93cnBrRokAf7vuvsLhEcsmw/vfzNJMht0UII/4EcmWnw3PZ4dcNfmGa/HG0SZOfcD43VUgModEZa
jm7w1BD7Suz/XNvQaKvFKyLwGfk0kUjcqQfq3gWht2/0IWtUyHT2rGhHUWj34PRKLnnM0ZCeDbD3
YV7jy5q9dVfffEFDrYsxXsFWMeOES5tCr+bh80j/GFk1tBmMq299dQu45CkL0ux+uDq9h6IbY4s3
A2tHajNodC3zR2c/8t0KxuuhHeBfD1OBhC5CdX1/Dp1oIKfcvKRKvvwN991Zdlp++Fbu72HXJnKq
IVFRCDrD0cdH+CNfi7/dpeCVImSgXyaojIQ/QKtdKll/hu1sFqA3TOF+QF0DNEK9GCjnXi0QvuWF
JOn02P+OUmYZT6pIk8iJcbF0yoQZ0D96pfs1F8L588eoI7C9VwYEnhxgSLbVrlEb6wfBRZiPN01x
R9wtF6wuQQrzWSt5VtpI/QjeeO3y4oXQmYgcHzZxW3w1Y8r+ThIQVlfuwCUo46Fj611a07ODiYrj
A/dsKETDb61QVYc7lBeDkxC09iZjbtVhMnzlYJ+8AN1pHMRkUqopUEcGHp7GtYackjEGtr+EGVD7
xztwb7cc72Alr5uRc7X9eIMdYdSlg3WmlUFjLrJFnAwk5eWKTOYaeuSm7LEtqszD5ZhA/LZN4t4O
aadxUQhWW54Uu//l6VeHrAa7AjvN9mPBHNzSCtkIoRE+rCexsvT7EBWxfE8nZnDr4xmTseAGg8KB
ciZpEGtXWglsLmobW9OqSZ/vl8m/PzgU09euP85mnK6fU7WFJBH/YtILWOsDKOb84zmlu4XnItcw
0zwo5K/GrZidjSxvuJ/DyM8cWCqPl0TQ6+mXLmNvr3rQedT7XLoUsBS87EwnD98Toyd1xd0jjayA
HjTVESxF/S7FBc0ce9NGYcvIu/0u1iLfehKUvbbiVDdKEDcZPn24tKXN7Zk/x4edNiKKyFC6tVzs
KOgCu9VkXKO2CRZHBaYNSlOIjFnNHLlycCsD/NUamKtFBMvA+HkLk68pWsk1U7p3AmFt4Z/aeu1m
ITVaPAtilxSCHjCa3eNavIrHqnhRBR9TwU1Pb77989CZAm1CU0cliPT5peiCLb5j4v7Kgf4+Pit6
tX6CHbbK42P//QjZXr1vIgBHiERdc2aW0p9a9sjpyLvsk6U/Uaw8Qb4ZsEMJG78WUd5xlrqij5SN
1EYF9R1mynFeyDjBdHuTh8M+V4armYE8mOMiruvtOdj9eKEN6LbmqP6ktDFNS7y+FScsDi3Uo3qu
YP3ND7CE7KKMxAqUEwVmRd34bLinyOY8IhYkTNO3rIuOJFUDkVF7N6dgLbQs725VbjUTyX41nK/F
pCBC6r/k4j3tJApyr8Q8pUd6kggGUlAn2elRmRsTqPFfaKmhou+ACYiIYcz2WMdyRtQPx5ZBMx5o
tIr/I8vFDIC9QS/OutAFvmmj5n2xidYNZ3xoqh5nsLAZa1qfIT+W/FgT2q5eaDRjhJnK/5R5excD
x/Nqor0Ga+yqVZ9jtaFx/jtORwfbgl/w/cnlnrwhf9RY9DZbkksAtlZY8yoPqtcyQtOFMoQijQzJ
9vCtDcmMLNJtPLSQZUhQHI5fz27ME2/hBn2Ci8k3hKtkl+/l8V4cs/RV4qEnFLBQKPZ+jmz18Em8
Xm6E9BmvpfYgKzTBrkWyRYRTmZaZXs3zbLIQTq6jO5DnwHvMC3PsKcGvH7OlDkKYr1zqGJra9QTt
/UReAuYsjDyCpTrmmOJ7xrGDL7qxxTfcQqWI6u8vV+lVpR1v4F5boIL8hWfscoMhyXG/+0wvSeLJ
a6bjeK91ntme9Xfok2FNWKyIBLG4nXW5+iJ4cjXe/GdLBkuar/SpOPbinFFP/Wk0ykyQhmro17sr
wS9csh7cPG/TtKj5grZUKUlW4z0MrIEAhmTDkYRwVfJIUZcXqAQqIdU1S45DwsPwqLMIqQomAI8d
uhf0Z7+R46Szt+zBqWI+8IW2xZvWJ3EWSZP3b2JANExqsYGnPp6bFKXLHKfyweI961lPuQXKNhR2
ovUjgHvSJEy0aYd8YMT9CVVUYzzOr0QkbQCiVSTsrF1h7jQPP9jmeg/ft5X7q+8ykStd6QL/rkxz
mCxaZAvIJxHu0Ex+xMjyvz0Z063p9EFgm/Zn7n2+rk8n4U7UELjNwNolGEKhBmkEi6pBtRdePdqL
NK1pBdPo75SrbKqx7gcLnBaUHvKDYLtu25d+6gYi22+jGVH/9c0+e8h667DzXJE8gCwDUUOR3GAs
OjUjYXnJuaXuV6D5iKVirm2JEEpz5INltITuW/dm/nM385Ws9Fj9bxyP7gspa82+z6pORvGFONa5
mKFAzBZNYKE8wCawost8QSRD5/zX2qPqNBI5Xef6tyQd7zuzSlwzCyT+SbWMCt8T/q9QF09gft8d
KCoL93KbNQ5sQKS3tUc+lW7CI2KdzJkaSbSsdT29e/BKOidV84x/Z78Ou02KuEZqy+8Tmk7hmgOB
7zweHqE6LVqxfZ1kjmCdksgoam+yz+NZEIdi6lc5oUYMptdpiPOxDXKSEhxFkaD1PZXnfL6S82Bg
D3w32B67K4Cotput6zNLJ7WLrjnoxgY37UJahyMwx/Jw/29CV4lcuwN0+rouLqbzDr+3uJHikghA
RsWkKLV6RPXqnbyLKBi8MVVGogDGusOeapz4ALIxqsPJGVDtvObCmy/FNFgW+KcR+3SeEvmyWcCt
ExDd2H2DxFElw355M9gKRiHWItMK4PibvKj+YtYsA5OcVMQ+nJ+qo4a07KTf3zKSDEug9egFxg0E
a77QQ9KxbQVYR2XSaO3RXpkgdaxOlWjhnnVeWF/Kntt5APlbYO3IE05bSJyv3luctYAG3RMnXvQs
MsC2RIy66rquHe0VDB7pTgkxkqtcqhoEiHnW30pNKM10Iq5ABg4L+985dyn1ZqAZ4GifEAXA9mgw
lmtRyIzBVTY2SwDSqRXbyO0Vumb/eRUEqWZZMwzc0n4nkb1KXTFKhgCeecjaw6VijiJUlR1js2cA
/Emw7BasRSwBkFSBUHDZHPkiKw3GDtWvEOz8IfgoKA+57ShKBmZSpQgZqjVrCT98bdJDqiEg4eW6
my0CNrUdaaKskaXAnJ+oRHS28ZJdKwleP7O+RPyKZPA+/IMkMVf1jnBOubUCUA8U4j1KmZKYgN0u
dT9Vsaolgjr9xbgSL2isZobcmdsQ4rK2M+28+SG+Nj7xxiq8HwSU3w3Yu8WTQgqgB4Hz8eutkPDD
ephFugONpyo13skQQVrIi3StGFt4foc4xAfuLbP8GWl6N3mzGZAe5XUfiuEfGmfCMRNtbLPUPe7e
Y985NViyVTFRa9xVM3sQEjgNIMYvfWPldW342+lZ/ryzgYIkBRhH8a9lH/BQTzKIav9L9g5lWYsS
OnQY3cqRjokcXtGCc5xtcSxazn/F+LlHjzU9Ez09hK79QIVJEaTCqmYXDCKYR2iJg+IZ+k7NGZrJ
T3dgvuJ1GxYDysBX6nOSBWTqXaaWaw3RGG0mTXOwGGuxWlXRCyLdAfNwJak7NsQiqv5L3hxNhiGd
L4y2EGHbFDGAzU4HwaFJp4LvgCAnDsesq/u0EW9UWicXwFtj0EV6RHH76/l9LO1UlHPda7SBJi/u
2VcSQYRmQIlCoYssP5XECbVgIzLTjgDRuK8avXtOkb/dCxS2SqIfojMg1w46ywKQq+16bHgWEPd7
0Gh9bNvthSOU9Q8tuOJvi36pj1aiKNNlur9tRWCMnxK6J0UrYuJNBNtuOhIKPmp4q8941S6VgAps
CR6D3HghAyEVYbuRENUyvxzybREMyIDzJZEvOl5u8APW1iPdJIvynXBOR+Kz8wX4CO6Y0m5WudhC
Nsr1ZJz1pN2B7aMxzYlTIf8l3Pf59yQRjEgWrWq34YMQFa4KrBrHOAJu5gf1wbbryql7GYUxpXhX
EsxeCQMFp4/SZsGViRM8cKGihrYod9uEWBnDIv0gL+xvmUmPr2oo1c+zqVjLpY2WrO4SgHjg/xOE
CCusmfsjK7T+ODuanH1tyn3bpt45mikVRyUTZD3irxUkE9iGrjnK+6XVUMQTrtLKo/q5Thbam9lC
jBYZtLLNaSO3Pm0MArPG6vgUwZvAHnqXJsH2RunbvRWeYBm8nfJStGVOE0YBIvAHyo8mv2/1Xnzv
BP+r7TO8SCXrwFPhRDalPAnrgVGbcD9p8kFR707AxzV3/goV3ecUJedpbD1bYJAM9eaejYf6njZv
F2GH7k2hYfMnIi/3Bi2FcMpDkG/QFVai0J1mgI96tTuBXZhzJ4V1mYUK9fdbS1XwY7tOm1ZPtP2m
HJmMWWcM11/d2FaukEzXUqlRlFwYygOgy5gIXkiZS+KgZfW3xwZtdmfVoE4YzQE9Rg0tIdtwCEob
vQB/NsHdu1n1sCvmfQz3Ied9anz3+WqdDUdMucFgGtIURFr148Kfni6zYO2exBJpdKXLxtZRzUlA
6LQ1RGzDUhiWOkx/lf3rObSu83HsEmceZP+P1YbqmvGYwL5kx5KS0gi/Am0lIOFpg5XHMaDLtpWE
REXe/m1eeI1344dCq2mfx5y7I1dO3tZmxTpy4lwzTSyU2Sg6+nFW0tiTucd7irv+mSNjcNKu19VP
IKgqmMapjVklIJixU0A8uqsPxg5JtIx1awjtEcRRfh7LAhqls7o+e2p7ad8VkXCgeuKKNQ846GxP
Z6Q+KoL8nXn50Kw2sH7ARXoCbD9DAKpDFJS+0zFozBPgO9d95FNyrK63/+WKD4kEUD4/zHJ2+wQS
A4n9DKmNjKdi9jFH0GKIiarRku0qBfl+9rbMAykAgOufNq+3cSyPgQ/DP1h6HkapSVGP9fO0tm7t
yWlDOIlAdgY+PLFK0XXR8RDEJiCBJjskSBavtXYc0Pxqe8nVopRpKuNZ97iOuSLJpwavBicaVFE4
oIWXPh5EDOmh1z2GFC2g38+W97FiyZxKxlQZ1EJ8WHdQlCVj6FSd2dBlR/uZaU5TRwox71oL5XxA
BokC897X7b34T76R7cDbjamSWoeV2SXouFQV/w7eUmA3wss46S+OJYrmPkDL/azuu3jHcrOn2OzV
aV4zhLXCFFeInnsw20IIggIp0tFVe3UU3vRd/b+3DThWFTJLxzCZq9nQsidFXzNQUD0G8MUi5eBU
KWCjLyf1MWlUDTdnZBCF7sEea5AggNRRV0q46u7OSodEoqP+s5Q4afpAmqBqG/xZsBKyjZ+kjGdP
6hJv9WumC/tjusNkG7I0Fc++DpFLfMwzueSx9pC5nLNSN4xwzCbAv5ovQcCQsIhnUOkhGjT+yLd7
ujlx0bzcKqBMeATGV6sSbQblfmWenLu89/NZj0ovszboiA7ivWCVn/gbLBe7XAxKZSZyx33yKyzM
97lFm7PrH2u41kf58yOpFvQ/+l26n+xK/fEG6a02rjfVetkf9ZfR39VTfHweRMyOlCIRGvX+JnXL
6WYUQl3xq6j6PGw8zTz2vqpjPxVVgd+OmKRS1LrQBhymQKlWNX7zM20mrVUR6nTeJuILFbuPByjO
G6UbU56CkuP+jTCnhWBpJ/LNwTVT41PStAe/vGNWloSeceoMm0IzCLDrYSbvudPuWWo0FTzJjx2y
9n85Kq9Bf6TXEmjJfbXl2spiu1+p0zR5JM7fwJtGai0xBNGTrwVG3th8b2Aurk3uJz4Ev+7kC/Rz
JbEaM8c25mveAUpdIvjioOCAeu1+wmtP+895hFrprgNXpj0Q+tKOBX7SjpsQYgzSEzfT9wSWSuZs
Ngf8GYTmv8rhJKf7QLl7Dw/wKRyom2WTw/TNrtARqJhTgsaVaT4hdXm3qoEJzfzaG7yBtfluRAPQ
TsImUJJhVNN4Usnan02yGyscO70GB+wLi3wjoHXMngWHc8AXJQbfj4dvrjm/zl0/Q57GoCUUcqZ/
29TYaZa/uV+vHQDrg4UzLSwaggHvdPelJ3fiL64DzX1yaQLeTRJQ1BzD4tdjVGhMHIrVcvnooKXH
Z11wh2n8mD1MKJmpmtJ4+yC7tqcXIqwaNp1rxQjVQVnCuF7HAKSBmHjmWvUmBfq4VjGQWO+pu6zR
YcuOKhj0mOHgF5kfPHDkuj8V7Mzsyva8Psiy/SMvgPwf+Xp8xRdvYoFj2yTndvqog+mlI1hVbkQm
YVIRwaxZksVmbxv1shXmezbr7O9+x1PfUrFUXzdQCJIFcrGdiVTQOQ31Kz3XBLyLDgj00NOj2Rrv
8VKixjD13lcRu2CWge8dfM82ah3LTWKDcs8LfnXKN4aTnZeN1kWAMXGq1HQPoEzFdIfPzrR/CxYr
xc6xlKP8t0XGKAv1fGi/8acJcaWdD59GdPXHJzIjoysuprYuZCIrnmcK3AI6QmFuBdIFI5YGonba
V7/8Uv5cdkwX6YNOEvIzo94x4o/4Zz0SUrKaWSnDDqG2odU6M2szNhE16Q8m0Tzm66aCrmEP9f34
DHQT7evuJMDlio701Tuup1vV1ApeEg7G5tr6Gg/u5ZyZVErd3EdS7x5Ef+vYbHsiqKfALqEGW9Ie
RHrrRn+qumMgpos4NdVx7p9+/VzSW7A3xsTpEa8rNsiA6QOYcspXTos3PL5zn3hT7KWoNOp9gAr+
6Eb6uLaBdW19ugi1+H97RR7Ij7vbRBCeg+P5l7zZZax5EgEGb5eJMteu98YaewtoIxH/v0N+N0ff
1TNyCyXLHJWFmyy+10UodSQFIetctvg0XrpGk6GecCgaxoBokoxp5ImBwxXdV4r+hg2Seaw7BqO4
0KT0jYXZ0ZKCWqIsp5eYrJnnlUPN0SokaX582HJWLA1cUKwgdfHMV5n/BRwg6YHxP3DnLfWQAqXe
uKvHnNnk3SnPm/vT1nTCd0IXstq3TuJV97cVEwa9EexfEPfptw0uzC7nj5Xf5mFW9IIURBGMF7vk
mSiYmXc2kY9feJvjGv7R2I8xV1mQZ01+Z8KGEaTm1y1yJDGOg7NNxzmmtFAMZu5xpqdzAVWzbvUK
SB4PXAM9SqMEwVs1MbQekb5pLLAb390SrP7RoI8FnEw0XVrA8dDOQLAEDUL2Ki12JnXU0LqWET0M
hz0qrpLUbsn2X8WmPPicL8pRWRncUfYVjuaQLXVRMc3jBPnKmz2BLVC80waEufeXJmHGrglcbKkX
k4pCjcJZE0Ail8riF9F7MKpzxXyD/m5SzNQ/yBDVpGqS4pxYdNaI8s7JxJxU7Qnt10VZn6K17OMI
pepf5K9vrwFT9sUjDJRUrywvaC8sxCaM3SZcPLUJCXScWSnTqunn1pRKNaKrNmKFxDwVYaA4uhxx
U6nf4jGxwlDzOFEmOSPqZhKMT7pVWmtfu611++q3TfyGfHQMTdkPsQtNd1C7pN0dJbTqM/DtOjjZ
qOgGtltRXBE3BOO+r6Nd/N3m+78rqd07M6/N7vr1JQ4p2IaEB+Xk4QrcuvlLgXHnsl43iKkZuFn+
1OBOQYPZ5boNzXBoOabP8IlFcuDipxQiiB6US9UX/L/2k8I0bPWooOwbWLEdHJBQouPbqxmzhhj6
y+R+D6H6hAiG1EN1zRJoU+VPxcgiLgK9+Nfh6xgfCmyeH3GhX+nwlwKjciO2OQH/DOT0yAdP6NAw
5Lr/oela0j+hvp6Z0/Ptfz5fGEzQDbCJR7zZ8dO91vJLz0Ie4NxEos1aM3n5oF8pvkQ12iQXESk7
iDHR7EWi4PQg5T4+YPB5vos5D3TFOkKfYN1XueAVASY5G4Q5rPtrY5/b5ap2ClOdMNHVNMzyzo+S
kvDAOFo9v7Ti9MVAjjwwtCqH/FifwKociVnEiiu0nQ9J5cPLcs9gGo5ADmPEfQab3z7QR1rE/H9w
npjDtibydw8TLxM8yLwTjApe9GGzQjENcfFX2sOpWx2VZTCSDTkcwmFOOq7hpOLBZKzdb4w9B7Nk
gNPfomfM5ic8dN9s/oN9OCLkbVA/RX1X5bMa7qf02XJq+D+NeYk1aRbpI4fD2pP8/fcyOZ3Rs3ch
XEx47MRBQaWzDrNyLr3jA85vaXy/nIbSlv4zVv2i5IqpCIE98xNqlBZ9/vYB4QkhgS/k78/Y7U/0
RSMYcIE7QeXoRile8BFg1vU2HaqCnyiMOEywvRukzCkDWDfqVVSVkWyfBsXuw38u6idxhUDQI89w
dyPGDQKuQ2Xvij6E/IrYIvVvCxHqV0jX7EAyuIBvKyhWdBaqxtO+fADSyijcmFynm3CjhMdaTo7p
5Atf4hXj/O5cWWZxBg3J/andTcDmx5k4HSPR+XnK6gF5Ey8pV/tOcPv+Q3i0FaseNZKKp0Qy0fNZ
Xxo7fn9zV44ypBN8hkxUFCKXI+iPN0wq2lGfIBJiZgDEUmqHLp6F0W6zGu9Vsb/d5/bgoT+Jo6es
eOo5w9FnYD8tRA8XRogzpVpFyZwEyje5+w/QekD4TZUb2ykcyMw4W0ZM4ythIyUUrv3sxcWcPIaR
dhisiEVJcXXG2R/pTrY792JPiKBtYFGPNbxQUSmYtWjiTvUMrJ4jBTmFP3ZCB7O++NgHMF509dQ7
9h+dnZ91j1SEx8q1xyyENdYd86IXRAIa5OMik6XoETQYTczGWUJrK/ku8450MOHfXiLZb/7HDhKY
0xMzLap7c49/SoeahC908ZpUCsIO5WNMiZRplx+Eo1HZ/ZZCRvp/pvmpcVqj2/QykGE/yEBiV8ng
Nn5GXCH3JHPtDFFtE562VN19f1rMFyTCMF9tGaWabLbrYz9+vl2S10L35gcHqTCu/1jKAsitM2sq
DnqFcS4wU5MNTecE4JtoloSmQbhpPdv/lyudMuIQV64JdauwT1HhRYbAbyJE/a2p2UEX8Hqv0Kim
NzvcplBtjlVf3gKaaZUSdBwej+frBjR4Brb+z6RrL/rG+R/DIW1DRtBD99XjRGH/6eFJsU49p0Tc
x4PvsF6kh1Gbf75KqoZpAkXG27ANHPdOfLIDWTk/yvbNY/Efp7NEuZxmz8uelkmGiknBf3VvamP6
d5OWontD/hE4uv1nD1SZZR2VlStctIUOTCBZxFl9gQcYgFGrbh5yYu1qfAWZ6gy0yiw4rH0APP3g
j6D0HmnQ8prVQEB8JtrNL9oyeIXCRPKrLA+mABEUzxdsITKp802cTOPKZUzjo7iv+QYbB4i/8MaW
oZN1J5fIBEA73cu5NixlnknjlCELTbh2BciEta4Mn2G0M6j9Z+HI8w8LAmLyrY1aFy+Tpw5Nhc6n
Falbo0dfvesd/gIrfEnOmfDTAywqDho4NM0cezhNjEiTUJbVT8umviSBk9NrTe0R5j8ZVyPz8IWw
z8IOTHA2SNTnWZQSOeoCzugFScSrl3/L2V8Zp+xliWdaGuO4n+Tj76AGR+wm2mkTAGDDnGSmLvtC
6NBaOEPUJJjwKrRpE6bxlBWNvsOv6mrocs3EnWvmNfG3OLLZWUXAxeNwSor+rBCmWUBt3UM5/plV
t6kXuW7bwvy+Fn0CbwKf1LjqoNs5Rc6jEe9RuL9+ph4JFdeZh8mBqVjusuxa9YqiM2RTnaNB16wL
Ord82L8OXvqjGuq07xJGkfz0qm7e+PGrpMPMNVX//6ee/ju6FYISl+HQiMLzwjNzWV0QAO0CRTHi
3WsXdWRuZ8dkm/wD3JPt+SNk7t//EQpzwjkLHaguoyhkOnuFMdg9YLaqzoi8mk1HFdMIsmxIEEMF
mMUsBZGyUVSUJiaV0cvMXL6VSh2zJHN2S2CO+FpZXSSF/FPxDZjWeK5vYS8QGjZIhrQ3H2xb5BU4
bvipNy2D3ITCyqE0JLaQdsdvpbmn0iX5fkyWsA2wP8hx06R6zfx2bP73Gci2mhPiGyFJ4E0L085i
cGnNuqTUfxLg9v7+j9Ji/RdeQlTonEDLmo0HTMXPZ3wnUJ1EG87WSJGPTqhJuaAtAfixLT4Ly5q8
I8/Qw8ZjKrhso/IHXhxWrPPlG4rNCjBTcJe4oWH/jlL5AQvNnUk6L+nX1GOxwQZbRmK5wSzQQ4Px
epj+8g2f0zvvC5x98lGk9djVERWROqhS3BVuaAqgX8xPtFOnLsbkUCKwO9T2TFbArHSJfd+M31Jh
sFUk9Oz+P1abO5ztK32z9hnhUFKIhPMUO111/SBVB7SbOd1a73RyfpWJhWppbSUJiQlPnw81tyVE
uo94WkpzVNUZQ5zUsh3eyaOsNvxIsU51vRJR2VPpdgexJ9Ek/l/fXrjxoN2Drwq7c8uRoLPuoQtb
CGeiAUAxWS+uISMvIyc0hY1Ff59y8J0y0blDRC5Gkdn+wT0h5vX3VH9ri6U+a9lKBWU7cmFBhi/E
2w9nmR1Y5wiZB3xqQdWNDeAqeWKVF+XaY7nO8hUsZOYAR2ry7k63yDYRGZNW6PkkcgO4dBS7Wgkn
oX8mo/vwrC8ADC/1/B9g9V6omLIxs5Mew/GDFULO/nQGKkVaIjZk8EzdVe5cM9dbBFiIFAkTTs6j
NUTn2q9he+ABl5pZ/rl6Orj3l5OvEpjTjEKDSWQG4+vIjOHcTb7YKjLh0KHbmL8IpS3mCE+kUskk
Eilr9V+yuf2lBE2WeMuTihpupPOaidXEmzWhLzzYgmOnG3b2+/jhQVXxwiKFpSvsf4E3z9g0YV0H
da4DQDbnaIke1leYUGe3vHueJJAI2ocYZ2xHPvBRAd/HZSsArOcGm6Gz43bIJvG1LLFcO3Wp1uM6
jXY6WpBNpGzSK/koR//H8QR9n2/j9rls+Uq3ggvyz7Tn3mInJ0OHOoQvTSBoI2AQ9mD6bW7l0mOm
A3OW4DJLdxFT7ySxcU4q2OUiRDHoRsU2/3yrZ9+L52gh61RMF+HRituvnX3X77Zt3xWJHAeJfqM6
ZMqK8qy+QkkhuK0vSoNf4y3kzEXzR1fJxuqBWkBUL8JFYcFwnISEqy+4Wz0R6o1q9S66Y2JfQkuJ
9+ErZZOAyaNQzdpTmOjJ+xkQHBYbNdwng0n4tCtOvY6eOUlGwjhU3PMir1+0jS++kaXThu9Y/gdK
7Iea1fwF2lLXDq78e4X/WmZaN7z8kjohEkeR280F/qDeUdYBGnev+JmiIjSa6/a21wZ4KjzfwnnZ
f8WNTERR0X0/96Gbj+waR2h5cJ3tTtzKgRBO+5KNQN2JRBxoamHgZ7MNBIQcRc60cMOSh195d1NR
thAk/GH7G0XDWmrvXRMXLfCvtUzWb0GlTYeSuKjKgQNDzYBKiVkhw3QaFr8hkVXPLTuBsRsrMu+/
YRNgi7Bkkb34aM0tAo7cnA+pgNM+C2TnbA8EJYgLqtKaXWZOCVtmSf8C+615Mn46YEeBocEo68SI
xRPqIuEIZGkhi5OU2txrRN5QMi9lrqldIAb+T9Hfb71lro55LU1Sa3bAYYTsjLmqzVY1RQrVaN/B
n1uH6BEypi5BVkjAsCIvdmYSwB8ksecI2iEWOEpQ+iDME8iSqQCgTatTZyU1j6O6Fz1v8TQ0Ulhv
j8q+pt7fpj87wRkS1dxpTaHda6sa1sl82ZfCAqlionV6jlmn1MyTyiiFp6MOL4j3o0pURMxHRCD1
EXZlgtuZGAPX463/aBMV2PzwJiMm+WzteZ3ML20ISHswSWVbHrpRJB7Jf0ORs2+RgDiBM0Y+UWeR
ylMJ/S+BSQmnbhsLPtq9M027dP29DHYZRmwTMimSaSndDTR9feUATavMVGHo0MtvWKmVIXi7S+Kg
hGYpoo0k9Yl9RIiqkabL2L2S5UKOQBPI2barRCZP/HIZgAxHvtqzFOTtwo0sSLCfYzOvxAeFrroQ
/g+JPvbnGNR8fwK3QjFyFWmAhTOovaZFs3L8aezw+5VtC8/mKUNxFDxwSR/l/AQdXNc3T8NSbLx9
/0cBWdAVII35yW698Cv4WMO9+wen+wF0tdTLfRKZjohkZi4/i+QePoeqGGBukDervyBhZPMBrV38
U5FTV11kyKM1th4vJyiqASZpTfb16dB1lkeCcSziulHkIVqTwhT160sAGCzlNFUk9xC4O/eq79Bj
V4LWUDBgqppqXIv234kPoUAuFx7pyhT8lhSNENLYXuiatQ4h1ZEr82UJpugDamGOdIZmxHBulmqQ
hspJWtfz4jBIb73J4IPHmGnoscwZuf1qM+LbgS2CmB4QjbaOSyHWfiocpjncp7uFB2SnJG/S0bSL
SwggWIuRquVaqrr1uWqIERh4qssOJLzEWUsGFTYTWBv8cpGRsUkQBxMD4mb0ucxZ95UdaMsDZDIx
oSUK0lRs8Z0cgw5G4Rmo/cvI1dOjtk0K4BUt5mpfRNjekhNmgMTZqJA0DvqKEp2S7UmoMuYau20G
UUve3i0l+xRsGb2gtgIsod7LYw+zY/pdcZUYTND2rNj4g6aJleXGfpDOTw56/e4nUXzJFBTcFcmG
j4wMbZRTqL0qhlE6L6VxBGEsXOeyqyPtLy6WhOD+R/N/VLH5nRs9bczOt+cJcrw3gwlDhhsjSE7Q
1aLJx1N4z9NFo8NbEVvQ0/VJK8FwqgIMUEcbcYVmVurTna6UUuI9eviX9XiwX5S0046fxPAjdWJE
Ntj1EK1ekJT0iwQWOmo+njf8WDWD3u0p2hMxPYr8yMhLU18XOb6OeCWjOynq7Nwo7ufGlbH7S+mu
O/kmnukjCD/U4BGTNvCUB2Y/oK3+1L44ib2DiC+QfaSN33EdmUrd7fVSLY6ST8HWKNccpdYs87GS
OjblIrI3eQXuPbAxHWztSbPa6HZkL6VjGedf2LYWZs5VqH9R5o2/5jIgFmqRH8msTBswtY83eOao
g7MUhct1q8gjx9I2981bLuqq52zOaZ0t+ZkVcctebjGj4Uh2wc1WEghVtUU9tC2BY3cIYAfY1YyA
xeAaL3bIFaKNlEBsCoJ4ZcaZGPWqr3Ew5Z8mmsZtvPAv3x3jigqxI8AQs5ZT1FsXYeo5w9A8bQJd
AIJh+nuKezynI0/Gl8dQtHNpwvCD08RnWL7eb1wzVIVcI7P19/thOVNmy26ud/xFPqJpCu5/Y/Cc
p3r2xfqFrlip5J/6MXJ1H/VBgt3QPTwDQ+bhmbiXHmPu4kJvRq9mVyfPHFx1Ob2KTQH01N57dMLX
bDg8oE2JgKt8EgvC2PSaDs/0EqC+8XUpo6bNNW4Cx1HxJrf6oLreJUiVx+O+tFuKjx3wkwlj1uN8
AFpJ9x9o0q0UzvvpHNCFe1s/IH2FU4Vy82lTZsxVM9JdTZUAj6o3Zz573z8t64VZxAUp8MnSqqgM
4Xzigb8lpzQ4ajlPEJFn2Djn8xDEcnI53YoHKz3/g3hxMP9c2o9qeMjFKVdCWE9Fb8E7qf1/daeb
6PFWOEe1zPKvLSnhLNZSRNoVvgfI6IYVbJTexczbJZ5U8rk6UPLMJ3H9En4AmstxzVd25QVR3ZMf
JtWf0OZu5A9WXgZUTfGA3UkucJXWb1KtifsjhOu5kEbjewaqVsFFn770sKt/DJsMRSdv88RZ2lH1
+zkr8LFbQb28It6PNbcwAKOOc/5NwBqOnTR9UK85QTzmOrmVB+8su0t5FV2PgMXRkqya0zUJb4nY
j/dsYOW6mKrxbrxOV2i3X6EE6ljz3q41ME47tTg/g28SlRANRacZ4kPjT4Ya4fvvdMK06N7wU94c
IdezfO8OzCmKqyrKTOFgm9MfEDxwCVavAvpZgVZ05yMWk2Ig/FDJmdDne52+MLZnTsy9k2IV82WT
Yo8+nJZ9I6XSJZ03iHY2FArCH2DCcVNUeCaEUP9HvkNGT1wDLJfHgNAsorHZJifSp67JoecKxPFl
DaPJbohp/U7YAq4nZFyRjEs5dAFJ2iDSezdFgsFHWRsTKJGpjMvYlYDN2DmChgC2IWbPs3DDWEpo
t2lneGILiQpVJzyoC/BdxpmpXyEw7b8bQxnkXG1kYACNPGEs8usLNLpySuiJMKZAInC1/4UTZoj/
MV8ihBpdDAoH8RI/qWkoRRzGqtnB38pMrSz2rv/ZGQ/vNUFkPH15BEZzMBSY/oE6IvMMjnB6uDsG
TV3YJIKCS2pyL8ru4VrabZx/exfvcwGGtvsC6P39y4Ja8ls3GvItfmk8qlvDREzwRNyVHJZl+79K
S0EsXDbbPEJX+0K3UZ4MPgOSR3pfPrcWj0KCz/J4ydpBgXQwaDBlE7eI1awQfoq2+6YaIq20gSYK
bJCfGjWFwwdhBPeDAq+JdnzCSsoMdLoI+u1X6IlQwtWDGs+r9NaXkWTpn4f8Fgck23VoX3KKKkNx
KEfaSWQweDzEvskbsAdL91ULJO1H1vrkbKqba2FBygztTLFx1n1DTHWuaV6jiKAK8D2mPGVQwS74
ZfBErJ1qd0yGi37XCiuh+8D6hztctquW2GLBULr2N4ah+xyGcNh+SCw=
`protect end_protected
