-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
cvMgi6UnJsjR5drZ7scQ+WAHjvau5JzlYzED1ciKn8PlRlLUdNmeti/CQ9t6kX9q35hVpM+yWBv9
F4xCysmwu4f3ixyUrusqrsjRqN7/70SriGDN/JIM1MDvIpiIqGOPvt91bQWaVUdFI2jR6QGttUvC
K+h7sRXMBjBv2tH6oHLN3ZbF7T5R3AlFtO0EKfR4joun27YxBPN3vSuOkwTNRBfOvzspqEeywIpY
wKtA4rXF3BqkBXFfjpgTmJvXikois1C1hqmDV6oSJMDcalf4xJEVzOrj18Ui1E+NrmrR0v2Z6KTK
XROvJpbYWxYRwyOV1Wo5hMjhblvNMbzp0LfDZw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5824)
`protect data_block
kuYx9oVduhErI3nmkwLJEPeyDe00hAsNspzBCDdkiOQMDt6jgeIXTV2oySjeHXEd8NwiBZ979y1Z
IaQ1LPbAiz2lGYSHwF+lvFBWkUG3ybBDqP+NHzeeg58ns/vR4sMS9o7jdAiRbDzZ/oiOoZTCCwt7
chWICKf8R5P3psLDC4dNpsqwVll4udwHgciVU/mscdDpdfQGJ6Bv53XtRRBLAYWbWiYlLBP/7Qep
5sf31+fr6QL0BG9FOoUbwb255jg8PaejTWPN/VWSIOkHxwro3I4igiHeHM5BhbAmq+dcuwUiRzt5
uc5rMIWAx8kISAhVjqJgogSt7C0IRBQz/2i28ZjgDQycU9gs1ZpR70fAT1yAuSjyH8jKWwbxM3dz
gHC4zvHZc10ydNELctEsJIJFqbLZ7oXzKNH+6BgSSlNNZXt5/zWQaAvHBEGSf8Z0JipuZ5RVTuJB
RDTq0H34D2JcwcNO4y9Dz2sZsC1MHGuOWBu6+tK2ccJZClE+nvA7p0W/hYo6BpwuHaUh4gWxhabs
568+LYlL0Eqx9+RJtm1gIgNaCzBOkVw6jvym5Di6rbVxGPe8FXPHzn7vdDwb2rUGcesx8yy3pBPE
6TS1oyw3JAWED8o6+AHmxlKZRJC8VjLMRRbIzcHo9sGlkCsiUxVJMjbnZFIh4FXB6buAgV6ScpmF
gaz3jrqURgA57meknsUdsKN+T/hZflmZ8fDLKb39H9tnfpNGrdLN3iVd3HSdJNsOXJ9ZJNuDpAwo
Yv3iwCpQJQoVsP9v711PDApe0m/NdNdZ27cuT3eiruPFldlIJ8jhP0oTvfOi/sf/vDGySqJIxaei
Kw7jqbZAYQFwOUfZtoRBvZ2zurxzq3Z+/r+u8amGXj3UdLFxyVqrLQe0gzPPhJeaFnHeF7QZ9TJZ
K3Z+HeYGkyupG2vDlRAuB8QHWiwojgX+VTp+08dsS5fSq6fIQa40d5Mkb9jsqM8sGbDYAoaN67It
UfWR4bOm8/qhbloo53IAJg0LWqWSUVGX3Osm5I8377XN7QpoWD3ZsWpQjT0sRYiyqeZSOyDbOKNV
X5mEn7MbaWgNI0zAd0/gFRBNoRSkXVtVkpMRcIXVUZE2NtnXXEieYXRmiNYJH1ekgd/PugMDlwxK
FRJnHt5WbjWy7N92gKYaLv5ZGPwipVqJ6TruKlQXAzVmgt2ljVVeYkngzP1spnADjDN34uWYtNw0
JstLBuIoOPkm/BfDtLrZBF2ObNSpqduyDORTVTfGI4pTjzxstPsdsRZ1zbFHvSMQXkuq9PCx7guB
0IEHhOK3HGvPGthN1rf5Hqn0R8wCzmZiYhG5vjyA09mCzG6DRFf6p3cByUm1ur3DMSonZYAvNE66
9ROP4OP6L3In7saoHhB99LM5Hf3gFcI4AeuubuZ7IS0wmcmYtYJi3/ovxBpb1Duog7sjCAJ5dZJ1
8b8F3JB8Xbigb+smuKGXR+fPsvBaRdY43bvJY4zhv8V20H61p1ctOGfl9zoxHA6vFZQaYLOYZfzJ
WghveEXunX6LvyO/IhE21oK2rMt974Sp3q/yDFpYYyyiqeN9XAs4JgvONqaKxGBPPtLRXK7g/lml
sEeulggtpHkcdBOAE9QhtcD78qZTGsYjrBsgpwyxkyH88AJIJnHg8wFpiFj0t70JMtPkKxqrCd86
KkcVpc1D9PeD1D92IMLBoPRcc0xvMM1q/SYUCJ7V0uBtNUPpGu2tCUBvxxiNXPTzSu0Lgq8bNseY
OZnR5dRPkl7D6AGJlD6rKaS/LDF7S4+fkuoJNza7Cdf3xxilZprS0NoSMc+qIrxUG1rjunCBzIPJ
gjXw9J+3XQuG7i8VKvU7iC+hs7PnUMPtyk4bVIV7BOG81r1E7bgnNaboZKM7kW6+18v0pE+BFiNE
wOu1mWfjH0Eoo5/j9+AgeXQ5vSpUXFw/TTsjwqbUqiyHz5EvMTxJtldrVdioFvKndbL53vTljXLC
UKU66qWSNUwkrLkEu4RmRdYNn4wPs5k3fzUPL2QyhhkKG8x4wKbrMQK4B9ZhPZ/w9cupEn1DJFK+
xdoKbLa31KUpMzvlyW/VXcClPMS8SjmpFiDD2HvdtbWLXcKSW3RqYNsEzhOElGKvhLTTKW3qW0YB
e6XSv9KL/BUi5EvX48BVfNYZ0cehB0OoAr3BBXgV/XK/JKn/h5xtOuvSt6gPlzzlWDLdCtp53zGh
e9qgi2Kdw+m7xRROKh2gE6P6CuPsh+Gcrjvo4hkE7uIuVgycTCNoXDkhiNpKPPE9blfs1DG00766
beDIww9THiLrelGUFtrhRp2vGJWN/TNQ06YurCR9AISqnSrgjvU0lZLgkoEq4pApw+dxGNG87AhE
9fiDTYFO7Eq/rTaypH2z12hDy4/AfsTQS8g6TH95n8iL6Jm58arwNXR/JbYoo3BhHTONvGsXyEN1
XsxxlrVL0m0Tv+seyUhgmW4nBIca33yoZCc2qRXBlRycb1A5/MCIDO0wuz9LgYRJHjtmfdW62+N1
yOD5svCW6LSN1aw2mPJyN9bHuQy7W1xsJYMVqS7VbZgwNOs78g0csgQ+ucwLfuGCmGQW0c+Ipp/w
ZM6W3v4FPq8F8H+v8CHe/lBJ0xtNTklbYZe19+8dgG3wQsafOXgmbmS+sQDhMsP4tbm5SKCz3Rmg
Mgnr8GcGINPgT+m2qHX98b2a4NUUXiZOH7HIDGaAFrjkPpPQ8ZepJb2fiiHzchPH6HgRfX3xxa+k
gsB2ZmQoiHgNP0D7cJ34M1MS3YhBiHOTcYnI2FqM6877qOd6yi9fBWTnuOwiK8VWdyHuWZBNsHUG
yzJ0q33vkLuiY7tCJK3gKlZR/kP6GRv0/jr8MyCQ3XpW7bMfcZRqUsYA2R1pNKXTDwTxSrrpmT4v
YqzCmVH3fC9CXMd9BQUm48Kd5gq1bsF57ydvebubV45RXhuTV8/Tf9jRSL+JoUaDjDTLBl/76Kim
6QG1+N8V2/6y/FOxZTi+JmQHAWyGzLPFcyYdpN0L8MHSQbooM+pM/r4mxleuMaYx23A+z0iT5Hsv
gzyi4BrYOvT1lnMKus+/n9f6AaIhgMb4qufhOhy++ksO6NLTwNaftmWC6H+PyFXMxMyUA92kq1Lc
FUAWqcmfTbGrcg9KxzoUadGoUNQhowvndBdwyVsG6ZpILLhF9WXoYv9S5KNg1plH5uHptqYtNEML
piRnOh1YLx37cj8PNLO4eTTZZnVH6e8X8tTa7HcPthC3bMDouJ4Cf8nk5Mzi11kWf4UrAeXN1vRm
6QszfLT2JY94cgv5Um7EgUHn1iPCs9buul/fL+mJMErVcMK21627Pg3I3xjaIfhJHlUVPem5y5f5
nMN6RO9+WhK0y+F3avMWo4YCnXI794D2J/mam4hSDJ+S3b19PNK0k598k+ZAkdyL+iHNnJPSQPQo
TM3guKaa406Ms6EYUJ6pFzZ/t0IcSlqfAqY5T7vjpaOcYOO7NtjDNeJ2APR98HbnpOtE+acE+8rS
tjEsJfDVRSoGnKatUh89ZiEXuPUi7Sa867/bs7vZ2wQVa3QzkU2gcwWlXL+Hq90LHbt10mjGDhfP
LWqIxORzFNR+Sm8jpQeaFxq720E+KKIRNNOeIm10jIbhEtk9IHNTOPsPqCtTyM+YzDgzpxL6S5O5
ysasDbqNMa7Hr4jHgSKQHuTUhhXo3Gx23HAAoVsP2K2crJzWrSccpEF0kzMh+bDGcpa80H7oi7fL
6eZat8zmr2x2OkZ1no+tgcF5/8EPaEptUy1QYAp1oo9JTaPOHBd/p202hnJ5dLcVCGOQaqypZ1Z1
3qmn3XeTmOtsiDgXrDK5xpHAuuxWHZWsOjYzICbihLCWR7Y3dJmy34UptqyXP1Q23mJfm1g8WXtd
BttsCiul3aZ4HWqJke19EQeAzWeg25ksL3vCF0ITp3GMZn++XVJaDTXAMNUTInsY6nEfR/aDIVho
zMK0VrFQyRq/c0a96NPMHBDuB66LnyzY3NwVuE5+zT23/okBnuLR1kZkX7LuENvzF46uZAlZGzpO
sWn1s0UFKmlhowmKVq0ZCLLCvEGLM03chccdo3xd2jh9aV9vdnD7bz/7E4WbnNjwuG3NKvUXg8vf
oCQR2u3k1Rr8jpTWBw6VdSk/tH5igaVxTErkozh3x4nAcaB1cnfkvhjxlzlNur8dREk5dwtVayiF
UyaQ1KKv6ir8PI6ZbRiXX7+4XBS6y3JQrCnQhhq5SzLTBUq7KHJVjt05EQZNrn64PKPLPSIkE0Jd
sJ61p5p0MXaS6h7TmOMCdwMR43FCjX8gI3viJH0sTjdAZJuTVBZNzQFxjLyb4tlGy+COR8Spu1Cd
h42CrYoB0XwA68L0bH20cIuHk/AhxWh8OyxW8Zv//OLe8aUQAv2RTvv3VhsjZAZM8yLzEq1zmq0e
g0Df6xDwxsmifyD9uq0oyHJKpjW6UIGBKGt9Qv1A2s8VVBEUvGMvgTaSydEC27ci/o7jWqOU5nyJ
JJA615RlcwNqfx3qxqDxOfchxuxO+cDzxoaDbJmUCqpLsvHkf/uJQXVxeZXyayP1qfgrfXX0E+RT
f7EarlDYn2DliAZZDLDB0bICET+weIeAejs6+3gan35y3UrV+b/F06l+J+T9XdC7zfTFxl5FjBg1
P4kE5Dto33/UAjuwsLFFP0IhgotetpN1e4H4b2oGhZbbjB12RVJBkvdi+AI0qZMaYfO15OyBhN0Q
KIpjKfBUdH2Hjlp2D+9QYfEyYMpo1RjXptCUxrEkibNLPG1c4CNYfqj5KrjCvQ3JAGiEyF+55GaY
TgoQp2c8E8wJarjDPbJ2ASV5KdnJiWXBjuPI6F4NN/a9gpJuSjDHN0UD8dMllBXuTTWtBYGYt/NJ
Cwi1KOiesG3JpF/icW0tGK29mGthlYZgnw5s+kKZQSDAXgyEgPhk8R3rUsplAlFfv4ZKSj+zAyPr
CxZ6hikez1Xf7EzJs8JoyOxumxnQLbpY0MrJwNjkwWN8lpSIeSscwiGJD58NP9KdlXr0b85/v39H
U88eBErh2r0sQF8BVi0HQQanepfanCr2rxMNentogXaGhsqzcY4JF2VuKxPfpZPm0MmV9MsUdTJH
kwHucJPHNx3j7J/77nbW9wUPoabbiSXp0gC2xZSZwnr6zmVsWd0Kt3kHDiyIcgo4MpTOMbmTk20g
aX8ucnh5/Bid8i4g2PHp0vieuBUJtjQnqqfMs3RxKUhHXZ7FAwVx1YCIVvaIhxaLdshL4JNduqt2
3gP77Uce6Wk5uef3Nfu5XQiQ4orHYRJvbnm2hYGwNtZTzODUQ2BgR29F/2huLPrJVdepR9Xm4U5h
3/mzmbPgX3WDsqVCxoDsr8dLgB9MHSWURraUvoDL06GJHL4RdvUxEw0F3kLSAE5eNAcvzsN6+yDR
PLMAoYS2/ZfHYlTB9QmXHIPbiw/9xoWTxW94YOA/AeOsAf8FLT1GWi3bdrjDq/oT0yAuJ5/F2kcw
dDgmkZZzfJ3xs1cMows0SqwBgELCSJl0c3P9XAtF6aE3xK6owR+1C+2gVfLCyj3tnE5qsQPWdBeO
wU4+k67xdEIrFJT9zrTYYlBY5HLk0wDWISAGiHAeL9YjjCpz09TQxM1FUtGMkvku5BU042A8sxHD
PAWBnwRhUiL2NGBctV6QTnjizKyPC0JfLZZCcOnjWajSEg8NlGrBNhZKlHd/IihpcKSN8n5NOuUy
+TNTkvQZjaIY5nPxWQE8oVilQWc2cL0x5CW+dPnnJpkYtogDc87JE8AfUkeFk2dWXFz8ZT5OpwHj
8bfHXj6qeqnOGCo6w81i8mPdT6acWp7E7HkyHagivFjjL99R4US6itIY0wEB0w6WVj3Xcf7HlQOp
5zaXQ0GqOWN1P/Z005RYiUqsw8CcZFLPyK0KyD1AEJKzsh/LKIJOlkEdJVs9b6jQDsXc54oZFt5i
zu98VgsQV8L5Pu3Y3jQY0hRRt5RydWkZBtVo4xoRiyC9+EHzo4zuwSkXeEPQ9uxgImJDdEBrSVGs
bb/d+5nYpKlLkpY8D/R0W6lKnzHC+Jdab2YtroqF74sm8oLa4cA6hWyzVX+rJjR0121YzYHfY0Yp
glh79cGGmmWXXJaW9TQl65OoPLfwcobagqe5F9/AreOtoMM3JlLdbGwPnHQo3wwhO+Qnk3cM45Y2
//X43KUjiiVaVowfl5ST6gDQADq51CfUZUmM0h8y8toMbUwYQNkhId5/w+Lr7Ixp4+iTJXkd1tXt
tajCBF4aoGxpsQhQ3HoQYPzjsPvVn6H0wXe9oAw63u6KPbVADUgpR6nMe2p6bb/d5jjUkR0ktlDy
VKoP8exEkxcCLjMNAcSUvLIBSALeHTCbQ1EsxtwrynYJWj3Jtvdkb0Eh9PEdPSvEWj1Dgfyi9Q3Y
F6DGRoil+Mprf1n4s96OH66/bFwGVeaHiUpgki+J5S36i4MaMpIAXwSbjUvKXLqPIzQhzbde9rzO
i/lpuK0MsHMVEYNzbNKCcPzGVcsilKTAMWHXCIDNDSqa0s405V685d1ffhNAYP1KD2SslzpRY3X+
CWNjPlEALDxGxuRfyR5LYmIY+k/1IS9kP6DJm8QgLvXSJq8e5ACl7RnH7lm/bg1gNCrJbM3zXG1D
kbzvE5bYgZHquWfbyj5EaO6ocNVQBYEv+DoJLtemb1ZLvIf8Fvpq6u3e8p2Gxl94eyxaHboHXzJJ
EnHHElWS5jzWB7sU+EF+hYGV0T6p93irCZh0W0JHBtlvFhEtsjoGMruXWtr/rhVkyEYXJCuZ8wF7
+OnkLrz73thAxZ1OINU0eLmallzsA0gSG/18rzNK0IvF9R9V/b/urtmgtS+LnPtDc+5QKf1C0dPc
CLDxnnurQCc3pCCtiROcyAOeihuCoymX3UyE2ThPiJxpheLDinIgNea+yREhgjbJD2jwSvBNGsJi
YCh4desI4mtEqTRvO/aL/b2heXZjHgeAvzbnlp6kA0fNn3U0vJvJiswbK5LiL0y7L5UDF2WNqaXw
4X8U1/otW2fxKswNes/oUJtFHhrVqj5ueXDXnMypa4SEg4CcuIVIR0/ATdEV1MgXBfpidWBQ0aVj
LosnjoWI2l+wF/sNSdLIf43m0yHlepw4T19DPDxy0+w9rc8oL6tclDbVcpAH2Pim1IwoBgFbkVBM
FkTrBfZUQ61kHRTdcJp3hA3MM45LD6oWNWjdkjsrng099VsLD5nQHSFz+ubQ4OEtNXPwSvahR5P1
8rCruo1Nz7NxF9UX6TAyfeVr5ok/b2OZrIWweEMaBaWvJNiriJeScmvAH0ppJIz9MVJJuC50VWU9
NdbF9soDMgnFeCYGTVD7uxnWx5+LyOMLyE9aL0BvG310vYbX1Ta6s8INxnaB6hZEl9Evmr95T2Om
x1WWGCu7cJxvkh+259rKXgdFo+1r5f6HJG80ZQ7fnOKI7ob08NOTmPNUa7qbWVWypw7dvdEcuLq4
Hb2b1AbfkGymEwaZQg0OLy20o0OeKMJhfaqqOgrbCgxtcse9HSmb19xoRe7lBaQGk20vFzRV5vUf
4kc2c880U7KGJyeZ5ZBJtSknpnXZPhWw4RAh+FpwKZ4ECeQ7J8ubsXeHHApJGnpHpO6gVjjisVt3
bQbP59nwjmh12K3he/ePBSN+LF213wxlypDT/uius1qp6/r1ASPt4gsf8GNxjXyxSU8qKroQ1dtY
FFgLiEYmkc9K9tQOVaSxgEOxY2RewWMstjWFNLH++A7Djspruqf99k/yG9sTF0E3ypC/BKJ5gyup
Dqu1bLxJbazOog==
`protect end_protected
