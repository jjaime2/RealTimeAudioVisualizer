-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fCGmRsMfEswBb5AttNpLapug+giTqsU0Aj+sWWCxxNptwKEImWyQ/Sy0bh2jajrZOthPZiXGGGNV
aYnIA5jhLI03zRWtmcwIeoV5rz1CDmCMu+EToVWbyL5KMJqwGLLn/85GVSOqLAXn5ooZhNyspB1B
WJNwTW4kSj9lJvfbOsYMtDSw5Fa7F/Q+YSj3ttweD+BngrnuVQAxR15x3CbcGYPzKuNSEqnSx3+Z
qXaQx2FRR7o+wS4IXwQdD9CJUhFr4TgUW0AdiG/J12CJHVQsH+3S0x4AScHOGpgeabUZv92za4kz
0nUHkVNol9digNLMoF0angcX5GFCjAZ+Nb7HBA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 49216)
`protect data_block
lXPj7Bfw+KJq+CAIjmwuXxHQJg9uegCRFk5vIRfyqxJy/xt+MsYXBa5VpmyGuw5/DIZQe01u4EK2
kB+V7j2uzOzBMqn/poUFWAtKeX8gUpEqQ1JYEdyAsm+ft0YtPlXfjgjGrDv2YVvus40+Q+OA+ln6
6UTR+EAQAMZywOjTk1EIVyyUhCB2OzUC85Z8yh/lwrl4jJggQaA7/MVn5AoQNKOvkuO0SHmNi5PV
fRubrpdlgECovg9Mxw0jpQQ1IoYDIWqIEd0iggkB1G7Usb94DoMQtH1sBEBIz3CRfz7hOiLVmd2w
kd+LoacLYobHOeI6TBazbr6wjyBy3HXlaBnjKtLP+rI5cmjzCzQLtT1GV8tAaMWuZ2lCggoaP0M0
HXrJTixDYFyYHxZGp9vAYzQ0KZENBpZQNAkWe9DwCAXDRZdpFs++NYT5kINg92N8OcvpU5VILGLG
MEMrXXMMpgrd2fz2qADTQPo6ptv3zG8mhpvV0tWkQNBa2eQfqihCRDuDQTJv36qzU8dxCOe0YxQi
XV4hAT3NGvhBFT0Q/wsJr0N3/k1FV8XeTR7oTyNrZYBhLQiusS2/5FIjRyTQLu6xDFL5WlUbnBoM
vHc5qYXSfwznO/R9/s4zAPy4YYhE2mbJH4l16xQm447SQ7KFq2Jm+lg6MnQpfuzjjloU1fgyBmLw
YbeTZTjysB1lrbiKUkRFUEadunYOY8g9hDJORPZKUcfgErEUBBSx71IGdU5QIOgpNr1qz7l2bBFA
1AJmiQ7aZzpU/VFNbzOnS3E+FNZOtDiA836kymeCItJOCGICA0OUAf+yq/TPLxYLxK94RlGXfHvi
WiaCtEsQ9xkV3R8/wQnFj8L6vgVmkaxGflx9aUK/o6RI26eT1snLsVsdt2aywfWQhbaKVDZVzlMZ
v18Dcl5OabLhnU6oYQLbzwo32Ud/kHQ/mP5ooD9q11EM+g1fZ1z7JcE1pGYmURTRol14Je8XlrYr
OT6d4nR/JBJSZH4lNXsbHTASkdvBUy6Lr0h+7LBNToRqqtO0Kenem40kQ0AAAe0cFrOorJS4eo41
GZTMG5sZkQyNkmXlMYVsgdt+iPaBuN2Kgq9+b0geoVARI/5omJH2GQG/zpHflt5qy0tBdzwRco9B
JuB2qDE6qe3zia/HAI2pSTSthrY7FUktNCGdCji7NSJgZmp7e2hIIhuxfwKckv1HaMDS0Bzv3HXb
qiFhxbMUWRgN9WBADeEm5j4FCYBPIY0XQV6B6FXlc71kbGkiiwU97LzeX08b2F/ja1CSielFeccB
7DhYVCn3BVQKMkywCiqtj2z/NFpFdqLC2MbHqFTBuxPQ12sg3ROmb42rijQvY0ZQuFj/9SeWOGyz
S1ML/w45oEn6M9srbx1v0VWggh87obPypqzDBh6lmzV8cKKmG3jBMiLsmtsY4NVHZMOajLbt/gi9
NRbqrN17XQx6f5G4e4s50DAMfieBDHmzp+cuZMOYdWuP4Km5R/GUI2L4dRMP7eiEyvVmITrNdKwa
oKi4JMdNdux3P9qCPdWSoV3YVIvxzjAq025TcZDnQIw3NZxXyVyXuly8qbH+XqPOezMrH1gJYJE4
uVQicCp4rcWdgwRDamEr1uoHzBaAGSn2kni27gGKf4VTvX5bALBTqDOteXAnXTGayOIDNLz8mFEi
iQ1Yl3HxWDJzLIO/jCIw3LWAzn9Sn4SgrHDMronktrf4IK/XWJNjRkmBh28edHHns543JTuliDLb
10zxT3B5RvKsycAtJNtCrW+tqJLIHbH9Vlf3y1Pyr2f2KOzOsZBvny0Ho/ViXNC43RMA0AbgLySU
QG+F2dRwhgUfoo4jIg9y1xBcvPyoPy2nyi1E7IrZmZsLXd94Ob6OBeALWEyom/z3s3Ocj0/YNKOc
lVFB6dA4MXiV5rzSHpYvrhLlNRCgo55Q+Y2hZJPtsvafbr3Ld54zuQOoi84PqVQu+YNNegZPY4Wv
z8gs9Kd3lxLlOUWTAJ9UoT3o0JTX2ZAvEOpJxZvQ6FStkg0HB10v2dmmgZ48USqt+R7klxsZz9Oj
t+EW/5HIL4MshekjbJEn/c/OG3weYa8DIfGrA/LIGF/VjmQ3ZF+JLjLeBRTRU3Krp+6l1UCnVEEX
GdI0sh4j1ilOEtmkXfWjrU5YG7cugXM6blxUChL5bHH5gRbHitSV0/BNOSevJQa/17hZdT3mMtYf
pPADnSF/ryztZ31Y3R3qTgDUtRvnnxwIWU1kFjKbPtgsvE54BapTrJv96zvtZjzyzF0H2p98Boiv
E7jQpBpC5Cw3b4aEZDPAg1PLd29uaWHLMEirAyY9XdrESnPpDWp/ttJYmZNZ+lYnYgS6bYEef/Rz
5H9n5POWbbClDrn74/ab8YZKkJueXtpnx/TGr/6no/HMZpcj1YDRzNtRAaIFuWErhfzOucLm3UAu
uqKEj8RoDEh/SnDQl0rauaw+4WYcdtOgWRazqkQMoLIl8Ao92pUAItuXNKAkqAc4PyPUAG2C85al
620KQfpeX2UynMvG1v6DzTi6LDM9N8aXmIGNKBHsROtnVboxVbQqooC6xJKGSoypwkugQSQJxmfC
/9i+8WZHYAWZF8Qgp50EadKZ3JdAygmjDzd7+37rl/kKDtr3DeR/lRQ6lz4vNNe1sWknZa++a1bz
zRci4LWtOvECquSUG3xtJPPjVOO7TVKvzLonGefbql3t1LaJG9ELQ3z5bHo09xgmq4c16JDOV80w
TPGDG5Zw7z/G9dAU8XnrkxIWtvnlnONLCqnPUHDBUMKLPFNH8Zkp0hFqf/6bSvmfLaYvdyztPQtw
3HJzDDwH1eUeLqOnt7Uy+8aYondYnAahcufjCupW4a2kG20F9F+ghkB1RZJI8kFH/H6OzpaHPdhg
EQuwfWT20VLutOpExRcINtazMbRitk6ABXYM/KFYYYjPCdCtYKEnWMUmvlQs77yyjvZCn4mGr9Dm
Uqs8zzPQxgZHM7Y+esDTpS3WuXprD8D9TzSAIYgnYjyzlOPWj0bLCuiYXLiOFplot4jWlfJ8yLiy
mQq5h9Y5HbSNinhoczbh6owBPRHAa+h3MO85SDCsZyZvwm0FHz0wV5nYAs8eLZeI2HV2M+XJekta
327az8fRAUYsNykOObX56IcBoih7frQ+wHADAxt9oDWxGQ6G7y0mhRvme+szVFlSTTzQiynXdO+h
5hmfP0hBlh24F60xM8Sv6Rz+vfUnluArFiq/xZb1lmKxTqdbIiycpsAE4XlwOKOP37DNyvvDb6Qn
CS3q+G2+PvqDiLCMl7H3EH8+qYlLOUvsmrbI6hdGCcWlqGX/GIZmL6K7st4oN4EPnxw9+x2762id
NV/XKTNAcc6W51264iwcQzpLl+2XLSS/yrleC26VaCC4bW/dzU6v0DENXedK0I4ofy6iF2MIjWKf
uft0/d50SD3S08/yFH721IFVPhmyupRjeNxXDfjreA3T+z1itNBgqB/m/iZhvcsNjkEsLh12d2iA
ySa1+Jmlz3pOJPEkArILGS6Da/mbklOTimQObqR0sZ481uxESD+kO8OySKz8nQEzM/nEnbwkKpuZ
fRFJn+O0wQhq7nC0NBTEtsbxy4SaJRDmw+CqWEAM4dVOnhsHy7GymgMCuOoB9HFCI7ajmYxjorO1
71K8kBUF/P8NMX2GZzdE2cXQmGOId24lngf9oQXst3ObYK1Pi1PptwH/w0fBRgyt9+uqWg9tIl2s
doa3+SmTaGm4Zn6zU1soovQEyAWo1f6vFlgAETqe29yBgxGbRLU0HVEtW4W3/NjhtnkrbifLt0F4
iK69SplHfVUfa8T0seq1wSaMwGzHoOLkfo+owrfe/rVcobn34zYVtOOoBx8Y1ort8IcNE6SAwInP
tksIt7cF2mxhXaGEYw7eX6VBvBJ/8/i1qZMKN4IkDw+iz12Vs/kOrrMlAuS8J+N2FU7pWqWqQy/F
Ws1TJs02pO0G5sDW65mHh2kyArbXa8i21ZLwgNzWnTN6ZyAgN3zYgSWLC3iJcu7mc0Vf8bW7UOiM
RDZBw9Nw0cFP0NA4aNBZk3f6vnAVVItqFVDk1JEihs+u3/gI7lcSOWs6A0AUpTu8pQ2SvVXRBf6F
PEpJ5EK616uPpJB9Q/jAtQLbqwpL3kGKYAAEYJC0LNBxLUL819ZFo/N7SJpcRs1GyZyq5i7W66Zo
hWKd8AvcKOe4oprEjk9IpaBNuM4P2UyVTm2B+jiVGPST8lNd69qsT7SBg6p6hKI/bfDvqs4hsSF8
HZhLGg9yh3xoYHem1fM/MwTx0ZCbjodbe9i7BcWHmw7xqpEw4bsr2pFDCqOTbZaEfleRyfeXA3gr
ZtWGqZwY58d+msWpxxYdC5VQXIuwfOuHxehy75b2fW50DCGIoOhwSOb80Y1MSgNf1TV7yyNwI/hX
/9yoO9AUPE2wxTfCYxkmicSCyj4llaCsmW7k/xWP3szlW6pcgWn1o50qVE2FsiS/nHw/8AjMZ5gd
nRhWBeBcBYKIslWNGqhOfLmc90TanUnPP/loYmHAvuqaTbGMuIbaF6/9I8BkGYA0Q3beHYGF/Icj
AeG+kRccZTZhkX5XdtBWTf5NjRRCiYt8lVZgsFjQPA1jm828sNGejgK3yratzhYuJ/CY6ipMZvPz
8by1Ld1M1TB7yAABp3ulxjCuzZm1Xhay4aqWvGy08UwvbgAkThr4y0rUFR9BUSpmOxZ14bQnPLx6
6tL3eAZ8SzjgBAV6Y8mhICzHNmsDewKPV17llxEmY9L0N7mzEQ575uAJNkv3z0yVfPjxALPP13EO
SDcOPVCE1LJZ8STxSg/UoP4+XGa3Tz5VNlfNFEJLXqUCju3V7U7jsM7UxmRrCd3ZnLtwmxV0OovG
yGBn0ZOC1hy1MlgXs80Zk0ZvalmYAlC/eMMpMvD2yU5yvJVZQy6PTz9dnqQ+fAz+ZdxnT4ntr0W9
uvPjxOi5TNIoplnTfrni0nAIZ5/3Fs45uhpFJ5vt4U6XrKqqmWFBpbZVZtNmeiwQOJl5aI4yjBVb
LCBs16cOMZ2V5jRom1mneqYPJiH8anMis5c6H2M0kPNFyMkuwJXKd1ovmQ/f7fJWNby5BjeD2EY5
8hRe3x3I4oYukcP6L6lfLG/ILtBLyuH0ndEczoMpf3hnmdDWadluQIPgp2zUmxrMhH3dA8aDecgu
VdbavEjy9SDJD0eV6ZSh7WCEYC8YLTESR07x1o4pDckz9zvkgbekiTuooC/uirh4E6hHyw+3Q6FP
5+Zg1kYHNfaHlQCdUOUB6yVKZz7/qAZGhuD/x073kBk/DuYc1cJ7T1WY3OEZCJNCdS7k7TkT4/gp
52+GNolHn3DZAL+ujSh3qZItRlvtsQEtBbBMgyFAj+YJefZ6cdiFculCQ+gXVqEFrRZQpzlWYyb2
hu3PElQBvv/Mp/MnLbMQmt437A+x9+rC3cr5JUa5hsy5IlX4RLedkBWVdV4dnFY/+nzEvygFEGC7
sIZQEdQ2tjw8cR3m9a/SsbBrVbjKjoNAOBGfUvJbkika0yoBz0jLuCALqjFOFzGJnGQoNp876mB1
0OoqOmXkT0mP3NRB2MQBl3g+XVAQ8oTcRBMplU6BA03pfnS4nmmI37lVJjufh9Uqu3uc5yilt3K1
eQaDvTCSeHAxGRBdHfg/gZktkrcn3w56w9lt7B0zhS9YmepaFgEd653WkUC66QAOc7xE1LQC99rz
/KDaBQwfkMOvWg8k5hUtqGQmn3yeuaCP/Ai6/UcEc9twR9LwzukBPf4MGokRQMn7OR0/8mndAZgX
FOQ57SUfhwZzzRO6O2lyw4RPP6/ovtAwxO+ZrFrgHco2IBp2C8PkXYNmIVHEThDTU171i5JxharW
DSGe/odPkv6i2oP6ulAVXYwKb2a4vhW0g1pMrGS1o6w9mV0D/qvCjGLW1UQfZSXLgy6C3HPmmctY
nZHDso5ttabiWmpl6a/wbaWFc8inXIBxfrraCVKLRiw8Lyp+RBlmPvxzb69k4CT6nRgu73mLuM66
2c6S7Yd2+l1t6KEQd7QVUcqY/WiapLeDghNSqZ56qgktqKu5qzG8hTCENuK+J/xY9Qp5QLYJmZLC
zROt6fIZHjNC1UFX2FUxBmNKFLd+yuECuCtFIub7oeeooJ4irtb0l1z+UMWrUR8ioT/g05QaHeof
LEhvHk0s8OA5DPbFldpRWR7OD340RU30ea8FSg6lgYGs4mwKJC65NyAWTKKtGuVlgewH5mTN1CeI
2NSMroN36I5tplP8gd+MbKvoMxS1bTR3J1r2JL8KPpYBKPyN5yDTp/oPkI32ezGzz+afTDBTI784
eJQic5wRp4UYaHQ3aVMGEIgqwJYu2MX8ClpYTH0F/tfm3e/+jW5aOdx6hy5OGUSh5DpcHvwmV2IM
zoDQ/T0cJvuZDD5lqvByMW6cNKSg2O0riOOpxKIkm409AJWAUpEvBHJvD9RfprB1LR+OSRMhks7C
rS/XJ4pQmmLIwKrtB3CPtULiDlq7wEwDMrldGRq5+niQKO+FrTTxzZHxV1ZMgDjI50LfxPl0vNoK
lLMuLR5GDA3qNtYkmmvZ+s5TjzgCeVZ2dbLDxXHQCIpvNrDRAbTY9SR9y3+kpnB2ajH+A22Cx+6M
7eQZOhwAMe4DrPg5X12y85SwGI1y928HQIICrhqxEyLxLtvgbhKR39g9jhpe50WXttdhzoMQ9WsG
3wb5KnY9ytxnFam1t7IiyVDiOV6MI4Y+yCoLkZK7kHBxIoxsYODtfEtyy40KrfwABzyNBH5xytCR
IkuccK82Qsls3fahCgkLMUChnyrhjuY8K+o/XP2lqDL17Zr7vHSaDleq45VozgUDDYkyZbc0mBDn
JMqKlpTXZTfY21N/KeTcj+8AqreVS7/4CtV4b61S6igCbNlpcHWBQCNrsYjJu0D0EvTW9jJDjd2q
40J4JxjK6H8z36zS71FW3zskYl+gnVGcuKbS0lgzVBWun4ns06J3TUhd8raZ87mRD1H1XTSj2OWA
yU75T67d3+wkTptcSgr6kQt8OS7HP1Lof6CrHrIR8EOW+m6w1lqPahZKKHnEo9Fn5XsPyZM4b9Rw
lKdYX0Db4iVDz0Wnue0uxnzgSMJNT5ctSBudSd+zWdMrU1lVhbA1oz6mzsQTsiKCn8TosKXZrVGZ
NUD7kNloBGX1NTqDHhU0rlimw7nZ9vsiKXvuOzZWCCthXl2BaghWbD9ahUmlY7N5wh9zoXrC0i3T
87IrxmhG5JkbZnHb+u4NL253wuLZjBcuWDfg8A4Ag9DzSa5lGXqgK4Rd80UDWY3XhavNdFsaK0Yz
bxcWtj+XU1OH0ekU2DCQtRpwCRl1SkEXU0oLcJSMBdOHcPFKv0Z/GobjJ/2tSrkMRg4uOLesbFTm
XBPaG2zb/DjdrCxWENNi54jvT1skkCqVVPLW8NSIU8KuCBJUpXhukjb8T5daC4+qB1IP8qEDwnpU
t84bZ1ODrbdHFcBNqubWvS9iyV+fzPygNUVSWX+YLe5qqqn/TY2yAjGVJ2v4VY0B7R+JqmVkmMjq
vi4oUsZCGjzzlA+Gthp/3wdu9+1WyvB9wtHCdNuYwctsOttYNxtLtfk1aEATZcHMos+N93RiRsZQ
VtXKMQwbjJDHVdjlH4UjThd9hvmpM4Inp6ttAak+6v50rlgqVb7FHvQ/cV1eQ9qZfIW+BNbQ6x4+
65mr1XgdkzAPSX8fUy0khagxO/+zUEvIXNWwucQcyl+OSy3qsFPTeKFy9TcIEaFLFgrCJX2B273f
1PQXTPN2+BMIY/AFLRTTRWqobodvtFm17OJlO0JGghBOpH2gM/D6P9saGDzSqdycok3yfrWrNp/I
V00kARR9rb7SEJKqG+SWrUdls4EddHuR3RyvUhmzgv+32r7O3sGCE2QLX8Rkbu7tvdTOcq2XUBXt
4xpB/ZVGNXsLWgLLpUii/kpZmVhDlQLddNCjxdvGcqRhfoGWbqcc+4hCRem9SzWf7KkaUwycDYhz
7ta9f7fDIwjgsByUP/nofybpEOuAZC5TSIBkv61/ocpgVDQnB0eIFjRcxmDvNZoTDYlM6dXAWKGG
IfHscb8zHMwrpuVgdlE/MwesYbqlSW4L9cDBycYDV5Eyy2OSGl8dV0xcpq+1hdj29zeqdTjJrKSa
qanytge45e25c3+rqwUfIZWKgwLkBj5zOQ0WqlfKECu1MXrfQL7Qd2xHxo/72KuCABZAi57EYmlr
dyVgEgIFAxzL1yR+fQr3U6886WZM8NmTpGokY19kdM8frVFtUCL1AnBm/fltmlMsLMYbv3A/EqSY
kjyOyIT06JbvTNwvN08pCV3e6tjJIXgmg4w9JhTUUSK9sjaUfJOGHM8c0upZaLNueUCXXSd7758V
cmCIzsvbZpcZcvlYnMf+g/Jstx9UuWHsKwEYG+gunLywfd5Tp/4yRJ9Q5wjyAmXW6PeU3FKGRLE6
bkf5/T08jiJmWPGautyx5dzLZLPgJsEJu0L26jqiXPy+cPGXjxX7t+VooSWjwuiDl42/FPblfiFZ
RiMu/09Qj0imwkNtNxJgappNprPrzMlvtZG/oW74drCerTjYn5U7arS4Osx7rc4DWzjnndboYQ5m
lCFHWHtQzfHBFeWov3hle81JfmWc7b5inzvvmT4/eOTY0aECeBiP5fMdPLDd7RZ/+zn1+NEts4LN
2iJ9N0aeaucA6rIzwfOi75iWlNKxq4DD4n1sPpaMeyo+Ygb+CYMIcbDYg0P/iL7udYm6m+L4Qm+S
yag+Z6SMxA85XuCcTa2w5vL3CLBz+CX7Bc5DEF75v06qXgFhNrsNcLpNUMgCkIQB3sf51f0E503I
Pdy2t9yMmnwGPu8bSEOoBfyW1Um8qTPx4tbWJS59m38yhDskAHGr/EoE2pM/CV1qbjuEUglqxalB
ela4cvfDTHFNbj3ujWbuRKW9CcsH95hERHw6CKld8nn6V51sKbe4/kYCqhdhji/8CZANVXKnuDtE
0XlGANVy5e3D9Dud5EDI4wWf1zG1+vUlwWSqomo4p57kWrM8523xxO6RKCazBaNIRyS4EWdG5Jh/
DXdd1/vpS7/5f6oWFLR5yDERjNjF57XKh+lFDL0Go9vq8cKvtT28yz7vvtDVvcHfIslwUcMQStMK
KWUSjgXEPTugo0K2IG4Yqw7jcLNCp+1C1pLerELZ+/30Uzm/zRNKm12dUWIgZgdOugdPYlGZ1qE1
Yok5e84WomaGzvAbycndM5ZHTHHygws7OToFXom1DOtIF3VgwlD1nsBXiJmEGvYhobc9LMQwTiOA
ZZVtlza5+CiFh5Gi20tWhbSWp1LuqesrptBRz0Slm7lsj/QK0ClprzLU7bc43cUy2php8l24wXt8
ssiSt6aybWJMLbqWun0gqhSzqwnH8NJjXliVsKpo7pZbo3YaDu6zwrfCaXr1W07F6/4Bd62yHLmL
IPWt08pIAB0LpGkYuexLopGNqstc/mS6tW+93bodb18CNJ9nJ1zirtygx/Rbdb6uQPkhT3XvRwCC
zmQU8wR64BV7QTdXa7mdH952yEtpRwl+iqEhir8ZxtCndI8Ms/N4E7DEJPiT7ocbQt8GOissmAuT
TOxUFHCPYndwwFRrsb3eSaX54boDYFyPjMNgcBXEy3vr8HJdbarFzUYf+HXNh0Cuhsjq8jRMruzu
+1rk8/tk9jp7bTgnmZ22tP+U5K6w/LlfRKT/9zmFOzzmUmmpb6Ux4xmaWfxZOGX9T26wnL+rxIu1
yJ8MRaPHd1Nu56S312Dpd5sCnsgVClLwWgWuehUsw7iElOiYzuIcf50kpJrdg1pxSZs9BmZsjDn7
xhG/nl1AsUBtYoY/Tf9DcTPFKzjjvngYyN7bH6bgjJNbVMNuwrOiuNoflGTpMWMGdGXWWXakwILf
diQR7B1xFfqWWHs2z4A4lM8vKnd+VZhOhVvOqi7t8RxmHugTQA5RC9qpPgFwJ7SVcS/krlDCHixS
nCwS1KGXSQJzYlaaDZdWcqh0A3ETRek+f6elckTq4nBh6HxjojlZSbp+cJLVfbCDXQj6rOlPbSiJ
FD41E+Rn9k2StaC1GccjfPwhIAn8vSowel6Y8mcSjVfAtHnobHDxulfSaBkgHCz8hoKVAaHT9ONO
rsi9N6kQk2/tJPTHqpQpSArRz+SYjdRiWZdS+pdhGjNjVWohqSjQnu3x+o0SPadpZC3XXVMjmR2i
16h+WUEOoGrJDK4gYnAF6dhVQHZrsB6+vQs8ZQ/CHh7bhKuLtQhLp8DIxGSY4jbs1iJg/4aa6N4u
JTsZKK2uQMxTphCSKkRWfMspMvVjV4461BG7JWdW4UNKSBMwJc0M2U6dexk/kMUnV4hf7rhnB394
xoxHIkw3MRrHy6JR+545dbDHMVDXCZceIHsRn8ruaawszLRx0Tpk/vgy3GlGYj9ybGXr1hBdjzIO
KRMWQqKQKVZ6NLr6C8E1lbes8iDYJWqvDultPfE3J2A9b6Tf076Y2Zf8IAbKEWL2NKqUoRU415s7
vrWnO03kkvhaCFw+8uoDi9aMvCcNw+jdW4SHkKeTk2yC5gW82oh4SY0+UvR3wjz+JfEI8ii2g6nJ
cSTIC6tQyfUZjCYBNkT5cJvVMpNGAUenW+WpiC1uQMTsU5ghLTwMGdzHoKT0O74GqB4jqJDOmb52
dPFaMvDxe1hDZ7afh88E1UAWo7XvXEjj5eqeMcycUncugaoQX4S5T/OOx2HQjlNQadC3zBjxdFxp
/pJb46iC1ofovq7PMyhPCZIcxDOTuev4OC3nYvqnWpr82T7s+VNBSpAEs8qIzbExrP1+ONAjCeD/
RPbDxWx9xzutHeyPYmgpevib3+/6ehQusOaEH1EKUrxHCXuw56vbmnBtZtqAwCWwxGJtpa74QJof
as8mk5AjS9YPCoQpSGgy09/IubPXzu8gMwSgHul58UByigH1Jl8OYy2jU/slWz/vkC83/jZNDjIU
WXH2JDNcX9bfHGXSZmKhqUoD0v8Qc0Bom+ccB5Q0bUp5/6UZr7WWu59v3ENvKI4GCxoUwuM1Euvo
/+hca+/Hxaw+kCMEJI3HcQ6rXDZ1C8GermnhYeb0lWCrRmhNdW3txGfhv6216H7lcv13v1NHWk6O
TzbPdKTsmqUUvdPR+OvdA6CualKpjwpOBmrF28UhPfYI4CxdZRzZ0g2Z8h7FK5soKkxBO7DFhqMt
7RFm8uiPhze3StVNrm/h4qcGxmqv19fmmgWmWNI8tsgKersZDR9DKiyJj6GNEySHUJWa5vCrJyZu
tiyIWeJa/qvvuxcb9wkX+2lmSwVhylrejQ0nxlVo7KsrKucJ3JCYerVUiq7mXBtLA9I3GKMyZrgA
X6sJVu/uu6CHhvTwPL+YpGltXUy57p+kHsMUoWa/OnEPkUnAOYfpnl4ZpGsQtxrhVo9Eg4c1ls0J
+YIw2H+g/Ime079PfGvdjBGbDxNJyimgxRVAU0sdOS9fA4TRojoOuSlHyT83YJnpbKLf32E0vuJk
nwvkwclaTfTH7AF7t1Dob5CZSFD9pE7CJjY29piG/YypBBusEqq/wIFFMiX2PL8Osrip2zcVhQTZ
HkNU84zP8W9BjOOyotueEGjJJTom7omSetpHOz6N88OnjZ0L0Y5096T4YHOX65FL2o/spoHKdC8u
P7B0S1y6ORD/uf/x1+9RK0O+1CNYi84Ycbv6QVWTZlG3n5Mo5Cak//p6x4yVO9mGJ/MEiaUlqkXe
2F1SlqDJLLgCmbVy4asm91J7xceAXZyrOD54Iv/yKnv58oqz5nYjntedp8XEKecjwgQgFiJaaab5
pox4c8bq+fTVXvPwwyKUSy6MGtDHckdm2lodflrPEF4GWM9mxeJCbvGMdTbxQgrXhImaBW6ELBzK
hjdEWLZGlj4pSbWW9IWFXSEhHuKd8kznT5oWiL67piRaoiwOdweLrLB2yttwZRuOz/kT0HemTlgk
xu/xQkhFHMRD7Z7aooywSA+ugkc3XMIvlSpXcZC+VPUMu4zDdVJjUaOvm24/ctG8hvdvlGRGQ7oH
8vCQKja0PDAeuFFZ9B87B06e0gELPhoRiPMgWsPNwy6cyj9VrMwG+5nUI0O1yp44kVwh1zhyHOz5
xDh43Umhdg6P+3bt0q3s+Yqxl58jbd3eRA3hSxOH02Q1tWL2cm3eW9344g5Lc7cc9Fk/pW8o4dEB
OwLssYYFH6xQM142aeCLUNjAAIFJQP+Zez+/VuUltHHI3jyE8vviN/KEAW3bfV9/2S57lMqao8x4
PzQNcKBBxGjdNcnQL92Iupw1qDg6X2hLtcvVLbAO3VaVacejEtI6k+Ln6uJ9OYqlN7cGhZmh0Dmd
XLF/qXK65BTQ+hQYOmaXKNZl9VwpBfzcAYEsCkGRn6I9f+KLqzEFfHf7je+M/tPNSigjG7y5mWlk
mbP7/aasfEh4oIflW4dKWk88xOtbZU1Iz/AGnP+dID4tFOAaj67e4bil4YjRF2lwSXYlJUXdcJYT
K/upKtcju+gHEo/WpNOWg5N8n3oaDEcd14Nd2cD6qRA9c3ob9cotJaEAiHJrgHyap8Vn1JG5AKxY
7tcZ+3S/7vDkrn5Moq1rn1fRdpjR7FoQ6KdXIw2b0VmtJH4x6jxIJYZTCXHCUCk3zNmBXA2l+q6A
hHPAskzJToInmgfLs1VN2hjuBZyBACCDAT62Rp3R/7Ow/65r1SRGA5ywfywSGS8dxO+F+a8cFKeT
hGLUMnTCF6dree8pjNuq7FgQs2h/62FBO1eMBY7icLgDvtLuod8AAUj0ayXVGBPZE/3rEw+OmvhY
LxvXP6ZLoUWeSoG9RHJ78a4X3oV4EroxEQeARnlpe76xT/8LeCRZh+cGb613KMkspaFTGJnJ6Pft
eZ9yOgPexR+O+dEHyiGpFMMJx+i2HzTxbGhscSqQxj/Y42V1eo0E/zyHFa6SO3wPVTBEJ8T5RJjc
K8i3eMGNrUeCDclWAty0KXbe+MKX1ALSql/7dqTsVOepMgzc2lI75MW+HLDtT4XLzIeZu1TpN4xp
G9GpWWferghwCxwAO84IhDxr7ZLsZH59QoCzTiv4mWUK2zI3/y+xq1f5eg0cFGLRiHuhNamdngt2
4lexfIa4F8qNhPz+VA3geEWkBBaV44T7FjBIqz5yE7Y9wKmzb7e+Envi5UBwJBKp5Gjscxi16xEf
fvkdY4AF6hmX+hZKjJiJwFL5g+cql0h/wMakiOtuu2Ppu2nyOlLwgKbCk9AjQqd5JJWG1A4nqseA
bFfhPchcrl61+JhNHHVs76QUQjKGIeGkedamNmNOEc5NKt307G8LsJx7xyqiXsKl46qktSnXnfm8
luWMbwLwXoBQgW0uc6o/gSe2gllyQhBIpXsMceiWjdlbLbZEgWvSRJxvC7AvR1AB9+5GdWwPUxu8
RrN9GZBELVYb4AjlYpakB+fgPhgEs10YCs16laRKfPlmg/37Kfj3utchq5LM2Iqf506/crG97BPP
Zzv1YLX7brNXoaNiP8GkZKmVj3ojP7u8qk/WUFGmtTjkNV4ahCktxAjkEDaUDEfwqQorq2S/38SP
4dQTO/LwL4YVhCqR4/jW3M9qWq4vgA8C96BDgXOLYg2IehB6mGagLsKBllmvlWwwUq6SphKTY4Ll
S9VSmlOLSwrYVvPoSSNpIaUM/nkPq3nbWpC4NNcy1Q+/BHH+3xvNUZSGKfMfLBKQk4tZ5YsfOHOu
0srdNhC3/70h6Td/jk5WvxB6WW+qJLc9Ocp8cu7RWSum35VSveejLY6E/uLGbm4YPG7SdZJj5YeZ
5hA1odi2pQ6PUeiLs28K6Dkt/v0MhyKIcjlMVovcOiq2qmPlBlFWD4lQN9ZLoRIc69SzJnoLscrE
bxbFhzJu+ZkKNnuq4fbFDrmFU5Ydn5ervjqAFHS6wulDwSQxgBBO5uHOf9Zy18FQVaYhfgKEKDZz
jp14CikBEdruozc9N5WrvAMir5ZJFsUWgwVmrFFBqbw7ZZFi/VjTyn3o+w7cISR1UxEJqZ3rLM3G
jx0yiUFSze9d7Yo4relja9EhL/kuaVzWYW6Ay1myTswLPEm4W54J6UG6tOKvXTGN0XnVqv3i0eDY
uralfidJg2r3C5YNFkSB8nli57XxBkTp5Timisut6oZcEVXEszgwzXZZY9iMCPXZ9RWMDHQXGGbE
K8lvSY7yDBGWiQEUZEHVDcevtTm8/L00RwwMT+SD9QTSzzOxfdicqzplOYb9O6R8J6fa+UKnk7Fj
c1G6+fgp5EG2U8Il8G9wGuXAyTvhhYUAZUAkYKoGHhIvvk7+Y0SvQY59POY15BIb1apNBgrLp0wt
U/s1rM7THo4Laq2GU2ljcPEzGhzMIx5vs/P9UGx8u5jegVeof5we3G1KrCsXUe4n6ODkQ0E6xocP
vhRyDqiVDAEXcqoPSXcmu1q/WdUK2bvlvqWfOT+3GaOPD0nn13+T+eaiGu233YNWx8sLrvuDtANK
y6sG0/B4BSW3FxI4zMZ6bQd4LLe1/2S1sGl9VxAuLInw6Rki04TlaZ2+XGzhoHvVg0q/RU7doYWI
Ae3kKSuqYYspguv0LU+SriwXnfSHtnoEYU7YL3maxpgoNpwm9nwjFSjpJhQegZw6bb+aBMxLDU1s
G6w8lPp8W1MpjoLAhydTHI6bDqKE7Tx0z+dNnHZlNO1qI/+JvAal0pp0BcaK3V8AwICMSLqPOioJ
xg2uWqR+GxHxhDg4FFEwIcEg9n/VjNFCncKDTHAsGiwlrQPkCaLqt081NyUd1cLnv6POruIcZGl1
+pfHHlsZ3cQDmLiNI9GLqTR5ebfVcyiJbO5+1hBfqycd8KhMLtgdCU3wXgwe/KZopqmytUrsMxk7
gDrlNOUmDUOYsh1HQazLEncjRVjirQpY4CTKI7U1v5ZS4Os0R8NCZUMBwL2GQ9VuajHWgYG+6q7F
ovxOCK6xzV3LcNiafbZjub06ZKI7h9ecxAsK5QTWMFEw36ZDOKlE0lXivD+jE74SvdmyRxq7NlSE
XKfR7H7bxJppjDQte0Pm51FaZnzAxJGVe0dJ+mPYzE0z4KvvBrUO9p2fesW40TwThsUTYdO6eUTe
NREGXABVpqOyWzYwvYAO9ipbGYKpm+ThmQBK/do7xVQJczNCnTmJVC7tstoyCpVMGfTlw5NIoe5x
rSr1uIC8SLGTY2SVSW/x5p5tFoA5xgAH2XJ8N91J9OYho3fMuCEGhP0KXP9Wv8K+6uwPAXyxtZif
5B5kWCa+y12CQZQwFTDSDHtHKkgYJcZuVJGrBMzT1t5cKLcrCg/lpKQDc62XM2Q7JEw3Byq/PP3w
4Farpa1LRQHq1Gvr4R6Mjap/I+kdgWpZVdzErRVvMPcT/qX09wlySIJk3Hiz0ZX+e+uIxP3E4r56
L8XuOB8xR8auHH6+78Nn4P1LCWPqCsBen7GjuoNj1+0xJ8lwGAAvkljGP+ZWmEyw4K7oEi9yeU71
4QU+UPxfPNiw9GGWrpU+mhU8xR5+GCzkWOYQ/6UK/HOvnyCcznB6mQFUT+4GuAwzQLtuU505Za51
OEKZzyr+oSLrXSA/5UMZjf5DbI6J3VXIr52N3sHGhn8QiRee2IK6BH0s9aggGLm0KKxaJFyTrt8b
mbVPwQ1j5DXO/3LmWCNNpBxO9RtX52OkOaMiALdiEq8fGa1GgTQ1oLgqQonPJAPY+2iqsn1t82v2
t2DdiAYIxAQZ3ML8MpAAhI1IbWkNLD+is1u1+PgVjnS1WX66i8M+FO7cj9jkdIcHZGT73hs5RlMS
qel09iOjNQXSuw2f1lXmqdOEFLP1ox4FQ6G6BGXWMRwMASxkwfrCbNhBa4dmlxMWe17NgTm5Wnao
iq4Jxqoak+lH3Y9V3Za18MJKcH51H0mEVO1ka+AHAy4i9QUMntmvoVs4s9rZFPyAeFAri/zdWiN6
rPueh5Xxq8wtnbJmqBwwNT072wKn+DaG0GTd9nFUcw4x/Hu0g3VBwJsscANf+yNmydlrZN6+jXOW
L0X1j5qB0B2wMPd/jgPhxfgOW88dXJD9PEFMr3nRpQrr9IlwxznmPlPjoL5yqeze1IZiYAhvlRAj
47aZ16C52Zen9b6Hfuf8ENP0/B/TN8q0/Sd/c9UMkKugEVKPVvpCSA6/3aLUfWfXVsLu8Nc36nZZ
zVmqtOTCHzmWSAskVwtZpyHKEujW6YAxfvaz+8YVSeXolvzcrks3qHt5H2Hh1yHy8QiqKPlfoj7Z
6KDsf1cwOsjhQE2MoT8UIgNOnqEXyhmPVBbncoQMZkvz+OkSJ2oiblZ0zuQe35F4CDgxfy+un0/K
cE/+F3tgW6ckKMGOmmvpU8iOjZSFq3qkKYGUmFpqWWsbMwHkaWi06e3zlXgPOkk6hvN2jr15ZuP4
yjjPGnbHFBLgXPpaQbSetgNpLLBrWc0OJCqWEsfUCp+ddURC05WZJZ08MkuOFNfmy+YKUUsHoHcV
+irQDUH/4BTAfPxqTAc1K4Zsf+jwJvu4sEv4+iCNa48sehDBW9k6TXs9yGpk2Xt5j4TIwrTbx4KQ
IIhzby5mQKZ6WZmY7PY9nm8BnSvEDOOOMhSsTN8It9iZUyaPT9Xmce3TkcrpQGMZ7ZIsPPzUUW4e
NoCrvNAf7qn75iUYoyDacRsD4XPq+wTayfBdRsJPMgQQ+S064bo7qT9QzA6BmogLx9aww67292TS
ANBNH2hezQXjdvGjXbMZAfG3vM7SY3rvIQ0Bk5cri13hrDOkiyRrgp1HdDoboj4LECEOX1+3n5go
CUnrolj26zX7u7cyycf+e9uRl76R8YFog4lD3jCGzi7BlOk7RmU0UKHBKLqURvFThiRIVUF5cnPi
Pxv/rYIYPMZmbIDQ5SlwnRtVAcllT5vjfkLaXfBhxJzbxPGYARc7CS44yFdrGINUzaGdSr8GtjCu
1f7wu9yWJRMOk4Xvcr8oNnXsQjY5jThw7jyfINAeua16o68x7LHPD/JOL9R/kaXwE0BTDO07Lbbp
xL1B4G9b5JLYVNXv/4L8PiA23lW8rL8f7eJYfa4+aZbArvyJI53BoHyOFkSnHqAe190mfGvMdu3t
PqVRCngPixVukVYmS7p1vDtnfEhtMQKxIoqnOxlOR2To9E9MAZNaAdrh1a5x7ezdxQQN4dw4pTpX
QySx5WZrFX5/cL1Rozwv9IN9I4xdFuc3BteHHA+bGIvOzT8F58kl3KFJ4R0CfFVkAK8EdgiRtOJp
on9bFR+eP92AX+noEvKYyfJWxIYEWmf0x5OZctBXGxm2bNlDkFXx9QJ2+/9smvXXAYd/NdqMwoWZ
JCF3MrSeMFmTwr9+xNwjvvBQvFSRDMRhtv8xljWoVd7T4NLmVjchJ7Pjwco/vJtn5/gLSA8JWmsT
AVE+YWMvurLPiWagFVpbfVfZ01P2CBc8aeGJ1Mjr6xg3sMlbexxww/0uabxAgb2T2wyPD7sIC/hb
DGePmqeknhc9OEXCiCJYO4E4nIQ5I0E5ZoXrhK5LkTDwh11tWHYZnWQnAJohfNXDHyR/6QC3lr9G
fz3uDnikJAYcbuhJcK3JGXt/K2z1O9kq3wO4dntRToEqfagmOLK6F6ok15CgTLcPJjjhfA7m6IzV
JoPv7atV+RfIaYPbuda91k1AZ40OvzdZgt6OO4f+KNDg65gEHwanSC39F/wISUSWfqcaXuxjNNQJ
DPJ20QQ/tQsgwph9OeSHU5UMvoFU0lBiWdkV+3fSX7+P4pjUzTl+aTYqzWvHMGJXDfcGBAwd+pOc
/o9MfgZ7xiH61mVeU7zCAOt8/jDA8WmDiuWZlWJ06VDzr+aq5Vrn0+bnn4txauAey5sXaB7SU86p
4gHuqHm9dCZR5DAehslAcVK8xzAePEFCSIVOjHYGOe2xYtp71ROxfRIxbBict7Z8OA4nV6lUHB5O
Sfr2RnAdVL320V8ZvXxWB7XnpdMLtI9DssL9GYxaW0M8EU8py2CH+ob8PhDUUrxSmTpMbv4L5IWE
LT0ZBWQdwbQ6hUXue/bTz5hD/f2TNkKg0cGCzzNQCYOfuBnJQKMVBxEPSP3p1jkI+vgEwc//Jl9A
PIOk5yhFVCBOy8lDrjqpnb+b1Af2RnLslwEnSEM2AZHXkAtGS+7XZzr8wePkzchvPbY+8kr7gRm2
aOtZnZsj0IpNGhV63IFLiQ/PcBVv5EQJdeU9h0pHX2xl11f7+PMJhs1CcDwjUiAFHQ3ihe6X/0zp
OwshzRwLgaoGQ/alb93x4hLxIw68FyN7LA6RfSTUBdF0c9OvXJfMI80VHgCxzTQK4KMg/AfvU785
DykBe6AvhFsviISzNsddm3Fmnm7tbK60H4z/f/pwCTszVOPIjyDeSCaC3xJl7FNMfoRWTVxx2CiL
3y6Vb5VWTVVgZ8rzq8Df6RcZqCVgr7tqfHoW+jBs1uC11OitagraGaMQSEvWhVCI2VTDp9H8oqor
COxIgdOcOFCNTH+uNSNKWJa+YWm3/M01aDqfT9FKBNTqz1CVbzVXuOEKQq0aCpy4BiaTTid6rU7J
GYA5hnLmjMni7o61Ev8t1m7oYf3+teEDbAu3IzU+VJm0D+h5j0O4zALsyntA9xLJ7C+Ns215bL0r
eQAZbNCQZM9aZklkOduxHLvoUhxswpxFrdj4Hep4llFQkgckFI1ft3f9OaRPsYfNJYGeLy6QGjEH
YZMlOkeGJfW612ZQT0OTrQiVHGLADP1TjA3GuOM0ReTI20iWo5+Lklekg3X4q72cADElMlH58jDZ
AFFqsSq0y8uZ1N2miR4vR1eVKZ67qLjARM5UFO3B87jqalX7SZ6v+pgAUGTza213ryQXNlCy6Iub
ZS+O0lpenzWNihqFhv0kYMPNFwxdxe8RmLnonUqfCrZPhBiXSsTjGUj9hY9UFQROidM2TRdzlcU2
OJYJoFArnDF7vClc/QkMM69vYaUPjep7ZsNqaM2uusHZlds6xT9vea2gZF6p1F0JF0Q0QWXBP2Ys
gxSLu1A6eJI2v7h+9VrnOW9VVa5GmOTFttZVrjkjG3abJ4mZR4Ncu6uCnyOwL0HyAOTGQvNBP5AS
TKnEiByhG8aLSHAKocc4tzzddnbmAHFWLj7bA0fc406f8vCgOe4CCjOYegJEXmCu8oLkIXQmjLfr
npuV2HKRp3Q1P1BxNWWRZnfAJMd7qs6qONYevUZe45mX8r2nXTi3zsbcjyGphkEo9Pk7ZFMM/X3L
RlVRqOQg906w9ZQxrFCyx5ZK07U6qUGZ9Rl5S2qu5BNRE3lUj0oZXB+ipqr1CgQdndodWthxf94a
/+TVQPsGh/hXfW/24Qzc/rCIB9sdLg1qdCo816RlidSu8RIGN0VzioT/ebL2SstEqQIe+bz4Zmc7
0Kmrz7cUFGcv674Q5voftosCZo0RgrQOA7/coAXyIsCkt691Y5IhzG7IxTMXjbpT8tHzEciJhVYC
ej7ftMq4gNZhSThfDP23HNpY86To5xIyZgEvwWBp19x1P61zDJUZw2fS3g5QBEWvINBx58ttI/r7
yLxLjJejJ3wtaxv/zQowvcW9r3l7IJy6XKqitTmmZmWEvL8dfBZDPH487cvpeOMa7P1EoNqZHTYS
pEdL00RCJBWl648rFvckJgPpndLfzu5EAROO3Oe1V0Y5wg7WoXUOoSn4jPxymDaVbiWgdd8J+8i8
3LiUNtKqWYVC2jt2u4e0wlQyGtjUXrty+t1kFIT+Ld4ElbYSm+NRfccOe8akfirrBQ83tMZCopif
gcunFOdpvyZUFseIiWgvg3NcNiu8XW5wc2IL29KdwdLC2gwQ6ZVlq13Ac2VV6XmjUo4jNjOL8dn1
9ymgww3ZLH1hCQqQQ5yUUA70D9soHOlcVhd/l5MDVYAS96CDkjb7+N9Kke2ffZ3EveYr5LufChxJ
/33wtgsUJ3Jd54xVw3BGChSnX8kWidvjxKjMKYTzDMnDk6So6/LmcIjEVEIzh4uQAuz1xSeRE6+x
D2ABfa8c4OvQbz5irY7N+3qtca89A1lzwKif4br9Ly4EQ1fM+meLOXsFR7YYcVwlJR6q0D/UpJd2
M3RtJGZNtLyLwpUEsJGCbowEXwG8/gdXaZE2vtZTw0H+FazOz15EqJxv6iBO5QD40W1qcN5SmnIc
KqFbXKHfDjEniBUDkv08uC2rzNYcEOVjjO3p5J3GILaZzxhfqNc71o/M9YxuKtiQ9JymUS2a2Jww
P4HRJT5UQTmVkdBFyJQqyD3H7yx+9mtU2PYKau9B8SR7E4Z32FEVXKhNa/mDLZKbwtZfujZjeVBb
PlWygyVSTjqdkb7BmN05b9KKldAH1p8OZZ43rjFG66u4Hl/eM+yfqUbJXUmTydEIH+jmc//8JLMv
kP6M6rOdWtFjAdxVaqoas69m7mAKxCNiro9DBv1UoRy1hEXWjajn06aY+asyhjKDMJd3QSpY+oOD
QG57E+h0OKLW17J6NNbsbBLuSWQHnw2aVs3ARSmE+nqh4TXqzMBVps1ZazhWjtODSgwXbBn6yJ0q
3gjCnO25ce+2z+g9RkSaXD4LHJAT+bTU/4rMg8glR7I5p9PRZOjCgjGsHYWS8jo+zwQPxxYQ/Sbo
8mtNVtEqNdcL9z6redG/s95uZ/YWOaK6tnls2zlA216BmWUhHXD5/84cvLzzQNk0ZuYI4TKBA/jm
uskbOKGtk68UMPFdMEmNff6EyoIzssDsGvVw6t2XD1Cy9bdyOXb6w8MWnrUHSsDrmE4eEQYhJluC
tn+6ldcNxR0Oev4yyAP42o9kOVzxFW7c31MzMg0CIecMeVcS5buPMHlpKoQh0epg6tsdF+OHHzxP
CI74ctZ5AQ5ZRKyIqVUkEvdxTzTvB+lGL30TcTVr8gFlyQ++QI9G8tBQa2tAkJoFF9vjV5h5+haK
3M5I0Q6wS3c5RvjsKD8BCCuElnXFttZ8UgkHoYBAfk/1uvVzG8l7xNc+QDSGj0dyk+3ZQ3Yu0vXv
SLHeg3T3s0fQqkQPf8t8bi77adwsncEohxGsU8dcm0SuQt6MWIar4ahyIW1oITZpnV79t2tu9uXq
GrEhHVziRg4F6kxmc/ziFoyW7kEIoL9wIUApzJAbXlbNEZG982r03Ouy+NrEr0aLCAzzlSZZ+Wem
37AJS6nHXuyq2BeaI6EulRrFR9KoVQS0nD9q37Pc8RrVAYdle05SIWXCDBDyKJfu6fXJIoacHxjg
iJ/USRBpNaf/hYTfei4u1gLWqTUik/lqsmPcFVJhFVfWhz1QDipUjAoNcIUdElvwEZs3ldAAncv1
PjEhXiczBY/75u8V2P5oRh0nfEc2fdnb1fXipGiisvIefvQjTBNOzLPdqDgh1tIZGA87kuj1q/+r
kbkEsMsIh6YpG3ddugtgpcSeVetqIGmVfG8Jo1kK9SDdr43r8r5Tri4SzpjFiw0W56VJCfqrJeo5
xCOWlyTB/x6oQcPqTrMX3b/axN2d5gbqIyZueDNsoxY5dzV/4hntkyRrL317rxmovGky35Yzb2j+
W7Z43UIA+XTNqffK2Y0oovhWF32b+vb7HW/FItqKaXiG0Pufs3J7BPKrtSe9kQy8Pgcq/GzvuQEe
5ziXg0+3zZ7P11V4Dgkj7CA0lUwDl2CZHSpulBwjKSN+HDe45bqpFQpGJZXvWrBxxwGJhPdTkwp+
iFhjRvRf7xxXlzo3wdf8CqSksemrnOaISDUEA5AnZl+huJzl6nhrweIG4kqyKkBUhztKCW6Tss7x
VT9hgyf2BLpFZ9kDki4BHBKs16RoVQasn+YfH/U0JlEBYN32uxz0pZVN3ghq0NaNRBiDtEBsu26S
T77Xe4vLr5l490OflXaGFuX58RuXTfywnXmoTLO4Gz2lyYcaUsZQj5ZJLLPoqLVLOM3wDolG0Lty
wKQOeNH2iQMcDwpCANEkIxOhR3vH3rOxL6ja2D1QWrWysUroW9fnskhpy2cOHL+MY0GAs+3dSsiD
/9Mw0MeWU+H6A3Sp/MWHvZPrhWBjWsvetZqZyqP3VThTO4V+gwYLU5691EWe1xqZ9j9XpBo0quR0
nXjs1w0rA/1BO59KzvCZkl4DBkemLRzOigZ4XnjCyBgHfQxWp4DUdEZ4I4TZbR2Np/Rlt1MaYL+p
dVQyomGXqh+srYBjNnVK8zv/EGlhqEDz3NHKaE7eaHK62KlddZDgBc8DiPs5XsDROKcw86anfgci
6nEJiVd7xUx+rdXuhqSDrzfFCKK0GQgySoLIN+woHzKOT8fGiTYcQUXGF/AUXHWt5VfnPxS3samo
674VbdYhTNEOV/AO23H+eVW6oAuOD0LRFoUDVdARxMANNUvoqhfQ8GllfcFXgDqCWnV62nB+s2gP
X96xZrYCGzA5Sm0my2Z1RwAk6rqDYMqZ5ajutFdOCqvB1FRkXGgiBRYt4LnlCIgW13MgVqVyatWz
FV6lLpXz/8YLaquhca5IOAOICO060ynyFhjtIyqK/ApnMMkQHWaA9n4DZWSgjAhZqb2iaERSAdxE
4DVPgxmbkwlJ7NNLmj3fpZgNF0AiGhRji+GJWWZmQOS0zEZ2ll/rMB8vZvMmNpL7WwTpkplR77r9
eKlu8+c2X8ypCr1R2tjIA5F4TmtDtLHpt8wcMM0uwqaCKKpAM592bw8RzrwU1yKa6kAcvyluxAC1
H8AdysGQha4PySKaA/+fNVKBFFb5e/z+s7LdCd1wTYNfxXkWGHoq18qG3kSVpX9nUAt/4InYX6RC
yRwiEagjvySNg1aovnqYfZFI0OVeYWC3isxbNutCMfKyYyw4up+OsSde6rIw+lkGxhNfUSNYlSZ2
PXAtEFXWEJNf5RpcRBTIL9J8XwLz6QiNVNEXRMvl/O6Vtw0AKDxRTp1uJ8SVKFIOtv5L8THNSR4b
KyBiYXLM1d67S8GwCSKRs/Et0EMMiWX7ceA+NShhsWFK3teZkNKdymEMmOkEr5URo/lmenKU1Qed
Ai7z9C1HPMx2mk+tEo53Stn7DXJa86J/WcfzrIVC5rClA5poc2yLmrZW6xhz42ryH0rBqy/sFP3g
wWeDcKZ/a6w7G2UwcT4WvblRWayTRrHncJrly+1pfqh2lgLqs/qk7x/gDfo5crXCmiWN9lFSxEty
R3FPBRTrlKUydZGJ8MjTkhTaY0gVBMdp0k377O4RRQiFUazECHQbe0igOGFeiGfodSl0dx9oiEQT
yUMX6A2/gkNhSbTNx81BBCTqLoJXzA5KeiF/3sPWL11TGMQvPI8SM8q4xMlcfn4x0r8NNn36EFze
N2CK1vfZw/x9SqbH+x66/qo8aILpfDD+eI8nqhDr4BBNC4x+uCtn3GdBHX1+Vk9aRxD9/rat473H
MVlQMBjBN0ZokpTSPltUnXknxbBt9dUgH9RQb0N25d9PbK9BgBeGELSXxZ6+jQrDNlLm0PZ/aoHo
SU90lO5UcjubmY6rwHQk40kILg8r5r7rxyj4QFJunwitaC+bEEcR8bT5N6SZpKCAiahbKLJ09Xb6
3eMOcVHBwUs7lO+619+2+EQyQxmtCes6ngyg7+F23FJr66edYbfJHRWiB3htPCtDVR+82xwIhRab
tCoxgI9bdaByZT6pdMwHYTHDmeicfJTqP24X2sCY97CZ0p6hNAf1JUdcKKsRv7PJ7IXACKGrpcSd
AWzlI5T2yYV83EiAUwSOatDP4ry3UbkQHdgnIs6lqw1TEpCxJvLYm2plJ2+QK+4nfQLY8ZtfxPky
dF+3hga965YXlQP1S7j2UWocwob+eli4yu1HAVymvRKIXRyco4DZN0pVZCyqRnLHI2R+jQ052i8/
aJMw77JlM5BrJXVdsbCpyIsEaMAF1ljxWqEiSBOPqwUfxYYg8OjFcoU6uzlVv30K6jtIJSH3Sg0h
qk0m3iXs1mRwI5INjWexh0KckRRa0ZZI3/uxbfulR/nhe9IlboQ0jnFCU9lGmpmyYm278ivf3TKS
ExWQUMZZz9vsYoBEsCbuTHndhwf/iGzdh+tN33Wm8XlD5lJcaUjbXy3dmwYKKq6zbd5HRhD4F2X0
BGGqArBHWjjFDBmTMeyRPuNXkDrS7+7lsvtrkSKDgBlGH93QxWDrJzuk6O9bgR3OvWqILuWMKDMo
xF+IUUrdTSZQINbpF+/ny8BMutQhw0lBmqt0CoKzIjsctvcOljAoPKxe8uD3SjbZ+BD9W2/kzJ5G
jABOlHeOHewgWsFMl9A3wSkyDi0gw9Et8KjNKOOM4uUk/4lkbfqKioERo0fPPxj4svXSel18Epqa
IZhR+tv7pFU1f4C/uhiNClVqKHvXWNbtPzNmzpbsygXK60FVquzAH41ow+PcR1frwfhztfm5xns9
H4kYC2RwAh1MJYXD+oN/OhuFNfpV5KnmIxuoPy3lUyvY2qgyLd+EqxSf3fqrdf0Xt4VaRJHnueXW
o5JC9KB/ImYKPaDsIJBR2ynZ39rIiJIS1/hHG8s1f1mtHkqbUuZb5IJg2FoU1tZt3YpU/Ud1YTfh
GNY5v9AeXzPk3Nm0pZpxwxUchVL3FkCOlRfXsWdPTvlGDdA4FXJN9yree7rVJIgRFdqcGmDGewbX
Tnj65P7yIpTV5hw0orHLA9gshkyQLr9pOdrePQ8YQ8vcjnr8LOITTInGlfCPeKq7LJYSzfrI2Bod
lFxvcz6YiwQfkSV0yabcKE5mBUJYmfJUfyPFgyAyzvMwxJPq9CeYVOqEHaCElgwoLrqADf14dOnK
EhPLCzFXWGknajtEFXfDtYtU3HaOgoSR0xYDz90i8WAy/vz9rkzSbFvBte0uqKbKj7YSud0X3PvE
NY9gp0a4UY8/UGOqhUfcie/CUYiXM6nSTt48mt5MnX270Qy+r+A9RrFPZMzf9HJKcGLTG77kXjVy
pyb34KXRIXygClt10AZf8tgY5WLz5yi8FfZlGS7F1q8L8TuJLyKevJZoZFbSHiABZEBUukSQYRSq
GhsXENllcLNKYoO+E5uayKARacKoqTuQ/RQ4vjdt3eZzULMD7P0bp78HE41zulgGDG0N9uUD7nYH
6atPnncJ7jSuIemXQgAelYFNnvs6ZAASZ8uXFA9F5VOkZVYsCuTuRZ79Kp9liONkQP82h0gspHxU
hrii0pCPt36FF7nFONLw/8H2nrxhRc3K/T/Tk8NAe8WW8CrHGdgccJMuUMvxgvL/P/1PuBAzi2bd
7yAK96IvvXRdIx1YRWxkuUxMc5zfcErr47xcP018PiCmJoUZXYwlTGV+xEcL646JJXS8RBD7OJUG
pEc9dHBwoV8TAs4XVeWGQ7bgQWsS+bP5dPGvEx+UsENjY5knAyU1uTNeqGcW+jISkS2SCxHAaj8o
lm+qyH8wOR5KwyEHJlsXx7RubVeJNs/jMWGWG/EwXKOjPgayFy7G0ip3nfp6OLYN+KZNJu6Cs7K3
v8ZW7pjSl1AV05DoLgqfTny/MyZ6U6bYNRPTb1P+BO0WNbqzP685Bfgcj84b6SO29X1q1s9LRVP7
WswocO39Oapg9QV+Ns1E7PGzQ5LcmUhOyckUkncquBVCghohk6YC4vZNXRwLZjOd+dGMUkfJHUgT
Jcp7MFQBFBhVbWHJxOa6E6YMapRNy87g8adesCwhdsuQ6rlwGVM5+gFWGiFbLDnYNupoMPbXv5vk
3ICWNskGqNIQ6jveJOup17qpjC8hlqEUFfy6Dr8T9v1NnWU9D0GhAHGEp6bTG/TXt7NZXZdc4gj6
DBQgmzsacjeltMUpL9noJRLHJoTSCvldbrly656L45PiE/uErzXqSz+Qz8yey7vHZhRG3x/d5WRs
NNxUx6bo9Yas/7Tp3wN4GibWVM/nHj1yoZ6RDmM+gCqF3f4o/VI6xLSDfQCT4jNAINpgfItd257/
5M2b+4+rVNw5afJApj1mNJ2v+W3wb0Q+aBuPHrR0t5W2cxmsHHmTCgjqW3SbcXlxr/dzwUCRdHTq
SMVgtLT8rG+Ku7gPpm1/KL1jUu21RUueRAMgUmMe5VnmcVM8tarrwB1F8YSWmcxrFYopNSeNoB88
B83dDHCs5yfsRfM6YeeoFFtmsOPbSkSLG6PAle5w4iZPnPfvYN3BXtCD/8Ov/IIjL9+WNpwQYeuC
U9ORmB7nUzeu2DBsl75pNLJ8nYeUNS3hAMRnKieWQmlp9S/ulSm5nMUO3oyY7o7o4jH6d9hPHTn4
eVsWtIab5ETNKIjHxR3SqRGbLgg7mUleeBwiDUOaSbDMgarDdwepGWUXlFGR3e1aFCbvZqwz1ER5
8K5OyJpdKnSbvi18L2vhwCkRI4jvVPRW51U8mlKHXBaWjq1uo3JTdDtZSi7bw93oboSS/XsgfiuO
XRGjUVYn68D50aiDwbJ2KDHfDafY2jlgltyRZRQztlSgKmtsayAmDa+aazGKG0kJgr5YAGp46oWs
CrXt1tpOAH58Rkwsqn4MOVhrTx1FwxxmsBU3LAey0+/DeoCy+1YvUTzFJac3X6bt1wI7YHjWkqMI
OXhJt+kPdoOrhIlw1wgq0NarguN4sppvhE3h/uEyvyyWv8HS4c1WwOlXqq8BCoRjuRmcW99z4vwa
3WDxi1zofiyjEIrtjxtqXM26YLNERL6AbXt/ypNlStda74Eac7DF5VRbeAc3L5Z0cMH39v/sSPZy
hb60vSLvjaDnzQgBDqk4nyW6hYqkRBn6ytyMbqe/+ysCP4dD0oapBtlVPbf3sqYfcf3tIO2rNudB
qSf34KUQYu6X5/8Ly8hfkgvsNvcPJsFsr2AIsv0Rj1A2BlLW1BsBtK2m1ttO8qTweAWGmy53Xox/
4BrLKoLp5s8M9KV6e6Qscdf/ikqzBfDiXjROkDjfJveiNJm8QKr3crKu4ol/4XlIP/4MDnL9GB7g
j8R+ozowBRNUkLh8VPpfbp0v/p4LmKePIyhXpBX+DTGCoh24HCHy4zwMamJBcLBfVxTD9Kl9r6NR
ZZVya9k2ntxY2gHYlbkJOu5iWTvf4GrYDau67R7fx/cVFXoGgBzGGZEA1r84/NWPtjp8gXmhhbKK
Agp0b8wnj8qXukrYj+p0ZyKvms6A9YWveUSIFQmvXm0ua9qOeI2bt/gaLKXtpcJxExhbopUY/NrI
dGNVjkZgXl9qOcd3i/Bli/A42o81vJduKNHGWyzOgdk4Vg4hHGEas7C2YUZYZapALTQjokbOH3Ue
4FYGXBEVv8g1/iwZbvMH8ot8j7m+Aecvqk5K7TFKljAxvXglRO76jPyznZQ78wVurRQr+2H2xKUY
XZDHvgJvjoXdyIgdYtwvTsf9RbhU8f0QBFFedApJlaruOEpRWkVNrz1hWV5DMKTW4PpgjZa7Htgi
vjBSQn0QKiTTmtrMp2FmucITa1pZChr3eTkFr/HcTYxjqg4QolsEAl4bTYHSTiycQg9cE6Rlz8eD
/JuZD5oK13lq2ADRxN/2iW5WMNvf9yRGyO8Xp9WegYPsWj+3Vx9pFn2TLivpJKCPCsSN98vRCVey
DAjrWoWLPZYL+HYeW8EwRiJ0c6Iw2krl/ODMU69gmFtmvTKjrx8rEeXgto6WqGBMiDKZjedTSPAf
dlRDJ5WO4YcbMbzqowUsV+PLOSDG3G4ZODPPP0Mqx8IQg1Kb7esjM2s1jW010O2F9C3L5xJ8Z0Yf
n3Ap5xv+//lL3ErgM4oWG/o9StbPd4N53J5imDiTbov12K3u/yX5tpJAN2ReJZ9GcadR2b0ZDVYP
XAm19REfq5HJXzq1MJkzE6q1IpMhBJR+Qhib/2YWTiQXnjTFZd95HGpJ9Gn092FcA7cqA2egDtJB
87MQjDPPjtewIa+JCxrq8ujt45ELfCfy9OQdqnJ/ZJUQxTyMSHyRXKJQY2mCzAuH0jIYWUxUh0Ui
WS7l9379Al8Ed7JJfHwoat496RsCrf65y1CxsVBPMKFzmcBCJTUPmwPUhHFoGLUldHYmafi5dIlI
rsqcFpa9tJBzXWqw9kJR9PFvparKVnA/8kE7WGk0hHZ++guCz6xM0+lEnNMkgcPL9mLcKsougUU1
EL67+bAb7gJWwLQirYU4YL7Ah6msDirkQzQAq4fsVpYB82J/5n1Mu6OVbrAwns+qL5OAOSxmP/y1
0bxXhzxvzUW9QmHyMlRwmwxUMiEApTSZCfJMJtk6R0mclquZvN+GWqskc4PR65jahKxEYqpUCl7h
AVi+qTc3UlDovM7HEZh64rgrqcxn9p0SR9MJAEkAgsv2jRdzmHogKCBjRJKhEZr7QUy/APwZoxOp
oMtxA8/lR5d0eKbxq317FbWsUC7/8GGmP/GkJMdk1nxvlSB5XHULx3NvKGlRHKFwC16OtPV9uDt3
ZzxqMYAduADpCBmZ+CLj4m39xTK2F6OHQw+VFyw3ZcuZyCQJS8iDahkPOjumYTBHrE1hUQ7PA167
GubgTMA613R0rs1nIWVmU0O8bUMUN/wp7q/IYJj7/FqwUfMqfJa/TFQqhgTcl2gKH65Xy7dG4V5R
s6OZwUi0iTe8ioYuUPqcoDuMU2+acVBXc0TfHbt9hyl5jEnkNod/dNAD0DIAonXwvyzO8qYNd2u5
REiLFTCdQljyHuOF+gX2Q9eRMV2gRE9HnPUx7xwW3zXQ2kbU7FpfV8C7SZEz/xaNdfIySJwZL+ky
I+JdHTIi2JQTpozUta68JDQPUdhn8hBcm+VY6WCf6rPoJLDb63DTgqmg9hq872a6ePReaIVS5CmI
TboLUHSHgwU2N+wNvIxS3HfNM6kGkkaXu8jzVB9HBMKxuvTv6fGea6re//66C2ozSm84UmFmFc3q
sgFKs+beEwluTcoRNnXY3/oMz6IxtKXYU0ODnniGSIrkoV5D1KsI/hTcELWZ5pnKid37JO0P9nRq
yHuOHSVqGhRln2baWV6iq+ELE0e4lziICkII2KXdSCv8dSy2o9Rfav2fU7kp1Br2Ge0k+7r3Dnhg
zIoQI6hVVszD0nrPFD1im6n0kEyR4N1O5WWYYu8ht3nvFJOpYGrbUG1vcJdsMcMRoEJ0tsZdspa+
zXSpGRJCoGtJGOQIZET1sfzcLyLj9jBhD3Bz/52PZtuTWNM0w8Q4U0Vxr70SwxZoWbT0t64n1OSt
YT5AVmfH3s3G7bIiT2kmx0CIvo6sjWEv9CL7q1+LhqOZPRk9PHVEL/f+LOP4F/8IseWl5Xi5rQql
+qSHplzUlmliN2m2/vBJPKJA/EAeGDLRNNBhZI5U+QmS7Di/DGe8a336dfrH0JCSXFsw+fr7Savd
BkwQmk3j+p/7dBV0o6aiXMZZoNFjqLbl98/dc1vlGiKinqM6ISA1FxEUQLi33AdYdBTsM/6fj9JW
vpTUWuIep+4fQcnRYX7nZVLbAF4bSYPn//NOcnzr7MoX2Wcswtz3tbjTOIvIQ4EECq7xeiym6kav
iuTtdDjBWKuToEM29ovOE2bZAFl/NZlZ42y81LoMb/a9eykwWw64I0yjmkZ3Eo+ZR3zLnbzuVkuZ
W5i6zf+f1JJp+51PYCSySNXtAYKUygq/0rI2ZrzIhffjbOTtzA5bTU3ihVBYDTd9kWsopGtBEJIM
wM6f3u8wRbe/O8KkDFJqY2N0BzuFV2osm6IzXXXTthJl2FIssYkyowQ8Rd7B0tyMFZqPbXsQhLuL
WItgE9SqCxv/xIKNiCl+CAVxUXYwqGiIE6o2Ty2xoO5sbCdZR/X2jB3PD6D35g/CT7i6uFz/uTGN
qnkhu0qdfcaMXfGL/nEB6vLEfgdBdyc0sFtwIinopxjro+FLHh9ykyxwaU1xxuf+4pPfh6Yp7jAl
w36DWTpEhxr7AuE1+aZ5GtI/DQ2Dx8SEuRLkYcbjK0MHi3kacTgwAvWD4Kwx74bHI0Y71QPReKZG
8yNnpOo4+FB4HR4/y/BY+e2iFvF8HJLmh+MoPrK9BvonMc2AljFUC39O0hh86Y0GLJA4R32EZxnG
R37aAsptYc9jFvexcgPLd52kC0TyRgI8xJi5ojZ6w7woMpHvfCCDrdqfp4jYtmW5Qk0nOn9j3cpW
xc8j21CZ72lPJZuROicMDRNR5FZ3lPDXPfLinnFFIvTATATTQvMtGkMDy8RKs5CeMrzWmdZQpMWM
4gidojAO14nEKNYk4/uMoQM/7PsdTCcbtu2VQOKGOAhwq8GiTtaD1u5k/4C1kAKNylhIYcN+QWmZ
qlR1MGLqfmeB5cTHHMuN1HV3rCr8OBo3m0a4XeqXc/mNtnSpQe/dPlpNTLJ6tGpSeN84EMsPMGpc
hBmgvIDiCe+KW+VizeyhneUzeomEODNPBldZAMICvkM3GCUcMEnBKs71DfvZWFqRW5LYLlne9G1i
SY+zvpMbYPAaS+gcfQkM8O5AKjeSm8eeCOpERzubUWFH+ZS5aGOYikfIOzAFu4VZv4n0dvBGY7bP
hm0SM6j8lVUqo4vv/l/9p3p65/UovFF3fgE//J3wcOKnCCh+/4EJ6SHnsNSF/ijcG1Q2ymrUMddy
4gxHaV2k0GQ7PqchT6Ju3/DxOtMDDZDCzR8io0a9fxwoCv7aEqAJv+bSvzX+V1w4e50p83RJfbvl
M/CsxfzY/9yIh7w4QP8b7AJZdPhkIYXw+eC9JnXNAB6f1eae83boqGM0X+fjnzv5objq6cwMrPp+
eFSPIfOrx9CPvdSEovUOd7suW5oEySQNttPeCgvRw68wwSxLklRaMxFl0p8b5+I4vxw9tVHHB4Za
sBw6Hz3uv/LlzxV/kd/GeeQH3ZILMxrlw+ZWvfFhtlLjw2pvdbapgQRWiB/1Y/EJh0vQxgrg9RWZ
3xHLVg8meKR0/muXjvtcQwxrBdwWjPN/FYspG2Pm2+ODbH/BobNRAT8qmwsWRpPjU4U3XF9AT6Cb
E2LF8GEqO7LuwkHK6HbiVS78iz29DgZv34geTUCnJdVP02e95BZN7S4m8lF0NPxtNxAPKSx1F1nX
FgD8Omp9sV42OZT9PF6Jw72AXPdIh2UOb233bj+ISBVfGt+B53JRK/hX08tQbw++Rct8pYf+WwCI
+KgfDUylluMlQAzeEj7v8TR11Z9ry5K0V/loUqhlSYxXZKAthwFZPbiqV7vzUjXVHqF7TGqKUjLR
wNOtmyqLcAvhbQX69GVtqELuZ55lJjV4j0eNEssyEUs1MOGIvxgQob1hLOQrryeFEf+EM8jXX/xx
AlXr0s7nHs5iyFz8wrLoDCycOvMBk97IyfMDbiBCXtH8F1wimu8hyUOAPPG0Zdsr2YE9nRz62uhm
1eieet4zqQm8bDQZPpFpIIOgapjZXy7vKAWMIifFZmAiMFVreCO/f8VdL6nZnuM5N4Y4qnaxLnqT
FGuvUI+uvska1Xvpyjr/M9isOxSysSvCuzwI0fLnc/P14J2pcSNJsxjMIBfCE6xrsON+mPY9mhBZ
uHLdH0waAzUBnTdQzfInn1T2Lt2c9OhaofiBX0NDPFvibhcabKuMqIFALkAU58j42XHkKxh5FQeW
A+194l1WNnDpxmdx1NBkf13vKFKjkPtFgrA5dXtlp7ivNa3kO/Qen8N9fjyZMC2KC4CzCQ9iHkE6
0sldJto66PPLF3uEK9Au4Zx9Df7TrVzafCQcojCl1HI0JtDT7Uyuyp4aFdZYftYpF97AZRwShqIZ
kmtypUijwHbzbi4HgDfQn8EAxnICOU0VzHpO+kZFI/xPXyvzcdA0Eu00ax5VR7eVfATnv+2cyHdP
ohrhb9JGTkL4t53rud10rslr+AXRuGPkl2lG7Bg0cWaP4+JnVreLjQzh/j8jM7ptfZFrmGRhg18Q
uZs7TDbVeFbAZVhnMdqbYOQ5DRECcigvkItSg5JrXSdSVIsg94E2nNbuuwqSKdFNfXErnQP3Si2g
hwKmyvynBdRDLA0/5v1RaZ+daklWVv59JKVUdLwHykB038OQUMNf1eAYDRtIxMrCYkGvHRbASXTv
AxsBK69004j0UI7Vx1wUcy6qbo9HYCZYm7zBjVYJxByrAty5ajcdnewshh0iaA9dYro29xwCMct6
0nVR6d1+c61O+AhnFA8PXKHuftCBu516J2/wZidkRhLTInnQZz1B3/syvVWBwfZgSnUlL7robSI+
gfcAPC58aPPG4p4UvUUOcuLYJS1Gs4wVQU5G6b3/XP/7F8KXBkaPEkSF/KgxRp2FtJN7lLRMXjwF
gKbGM+nV2A9N2Ktlvt0d9InyIpr1hvAXHzRcAzQOnMktWQUR0VeP+4sER1jFGqQ+CWpN0gKLl3y3
aE0biE65p0QpE1U/v1QlS3wbtUS7cgfcRG8sGlOUHOPDho2dTU7NtjaYmVJjyS0tb+BquguHLi0O
7JPESsiolRMB85GsDP88v0w/icaB1NJUBEd5h5YHclIEGb3mjmt8YLoxPRWJDM7dyA2p2vvumlF8
KlKV2NM1mWwBvBtZ4lAl1MWwiz0stoAuKJmagxdYA1Md/qUZIk2dXrwcqt+7+rIael4eESu0CuU+
g3GWTbwKo4G4a0HMiD9Vx/lFErhz6eIT/eMYLyCBjm2Z4C2PSJHs9gXXxTQ3xVPqqkPt/SRmROuF
wvdjTNKa4bI1rTYqoThVBHbn8KSClyk23iGMtUmpJCpBqbac3qo6NlNVpbBn+bg4kS8hYhykGRe0
41Wanahgm/eDcGZywlLlvdYGcplohPMxNMDpk7EOWHWSt0/SNryxa1OQDIFSyuJ4wANJi+W7ZlI5
ht9D6rnlCFpI+1OcC4JE6cdr+zjqcz8aXgMp/62b6na8ETU3wJAnTHWRWajkEo0BK46yM+VLVm6W
we+PBS2VMgx8z/Rdb60RqM1G7VWi4kw62BSgyI2R7ILp3X/OViXOPvhxMLbnpI69wKXKNs4hYuQr
ZcdaNRQVqmYh4sg6bfOoaAmXmOGmLk0Xh7UEzlPocuZsR9H3yNHDeRilOkooacuRKFzZALhOOJr3
T9jiOXTvzp1WCwVaLE8aC3uN5Ko+gf+4OXKeC7EuHdPZvTgsr5/CVZTfb3JJiOmvWq3sY9suFybw
B+svyh4CkdtSDnGc3n12iyd78VQ7X2kE+GXeGFkpiiBM5V4Ot5mvlN3m5V8TEI7v0fuNQ1FPzJeB
Ch8MA25wuqD/fj7bYnzCliiYxatJkn2w9B1GPnWkKHBdj1c7D2Lnxw5SK8L8xWRb6KLc47flVXK2
5hFuBzaQvGYoDX52tcjjtNqt0/ho7GPhJFWlaKo5H8m3FBdKWB648uWdvh095l6icuklxk/v7TUx
UJ0+9YZ9o+qTKWJEZ7K9wmTaRlTyRVbVJ3c/kTQIKGwkckw22ieZUPkP/GayASntZ8PzD0kLPGPt
ZI/gsTKoc11d2qDjs6bdksOXOAKogE8Uz/UeLyvxG1mvUW9Vik3GDlV6iJqNS3ECbe8toTuuktZx
aZa07xxgFL4b6eR6eIp2wQS5kQZHjipn3NiJqremcsXZeA46szus7muizHKOPoEJlX9LJ/5CE9vl
66CKkyggSWZCpRQ+bknl27zSemTIyjayz/6lGENLcs5apEiVETDZ2lN20PhCzvedpL6K/3LWcSUo
ua1JrvUf/PBAiiJhmEmZTJcwK9niMQp4XE58PgahL+2WMYsDnEfFMLHvCO+3jsVmskftyEdQW1it
OYfePnIZxLBQkZFGR8C3HjHCX6pdB+j9V/DOwjCVEpzo3stPLXQrFpkCq3bWxeDTcSVC6M4rdMx8
tQ4q9D28pt8ZOI0X2kr9zDVWCVdDeN7WBgRAcyRUEJzHWoyTJPfNU8ZbAxp01pdZGx5tcpSsI2E1
+lx/hWQAP91jMVWkFD6asc340FCNSodTRTE2+7er3JkwnMjwUDQCdmg/+uTqbvXiqO+uxR/N7xRk
09IxlUpuAz2MHbbmsL/QhNn5TToycBezkCaCFr+LkmU87KOIvudaxwO0Hza5ePSFR547GODgMpSq
sTsDVMim+Tav8gevn8/XW/QdrUI3O+dTMgY6t9VHiBDE5RoWdMgA2Cd5LehWfiDqmwJVmuTnenQi
TJzDlOMrDifmjOsXHSEetjZxLDZUL0OE1JGfeE+GG32ungd8sC/I0RYFumHKAqqllGOqiBacxhOj
tPf+Fvwjo1TIOEPFLDmbSB3vBggZs2fQdtRms7wy7Rv38/ZY3I4F4JorXsx2BqEckK1Sndz4TMk8
U56+mJ/HAOtFZfOW2y5KZfTr3ry3JXmhqNvuBua3hl5+vJpKOv6DZrOww6oae05n65xItdcP3qdq
4lvRrKj7GFhIx87as2/LbhXG4OKoCbM3Md+CBtWhzbL9ouv9uzccLVlYbC1KZVvmJX2FCP1ERVOD
25vlpae7BQ0hBMnu8etdzg88GUlSyGXg/KN3VvYbEzQjrlLN/Qb/1fEL1UWSMhigUjC+wDGn9no9
R9kpJdWGUTndS+wbAUGCgGtf3/u0EtYaXYFJZdWRhMtjSsyjQ0/uJS8shyPByUZPSq3RBTyIK8IE
pxEqlMU5RAtNRw9ay2aMCA7+lc7i4jcKJYkLdkEKpi5pmNl7smnGzQI9kLId6Y9bVfy5sLijhwdI
IK1+3l//byistnO6S2VpEZ5yvJcfb3Iz28YJt2oqZ9siBiZyyUAio0OKqHcGMfDL1FCprUnM9ZSM
c/7zY4f3WdjajXpEc8Zyf6Z1FlGi5jVkSeORLZ4ImuW32h1RoonNDZuUh/ZQ3Jr5Gl6wwkPV6vLA
D1L6KdELVMtOqB+CfUjo7la8IjPK4je+ImnTpYH+3hGhlk6koLZ3+7V6qmH3kmqifQLxaC5zfb0/
LAA64DplNUv3Tc1G2/UTETYZNLdBPop2gDn5KaXR8bRNt4pVwwtySUNfh+ale4BebloamgwzyShE
xxygm+Tb0rs6m1D4mbE+nREvscpptgA9OmuvOaqdcm7KMBatmXp9wHK3Pl1CymOtWU6VMq93W/z0
bFt24TxbsCSl8H+WmXOtlSA1xCH8QhiLtOdMUI73PV9m+hWYiHEMkG2MCjViSMwP+71XQ2LISJy4
uww6imhCILw+IT/K0Tt/jzrVLLNZhIT6ErrT0qD9jbhWrPZWBszLObPj+q1Byc+8D41Naf0cmZhu
p311/BxV8M0bdJ0LtKbMYyfoyVN7un2lAQdCKg1abubtgxoKBruhI2C6NSRvTgBq98NZTdNEagTJ
Ah+GiyhxsOXvGy92eXiuZ/plxhuRCJpvUJZUUQEYIeEaUD9qPaogINIrjT/Nx+ufEisAzF4Cw701
irRNkd7aeTFKPU6D/Qp139y5caoabnDFa0pDce2c32dkCu1TTNtT8d/xY0DhUui409FhvIuW2aBy
9goQimFscnEv9vrW8m5oROUas/BKLujdp5RboPzKT0W57OvFNW+8aj/FdRQnSnJnKE1w+OoQU3Fn
OGTryc07TmgKpCPwYSTLew6WN/+k1e4EFEuPckgntZFG0OeLnR+Esn6+dzdTtIYSvFpR+JyWC596
hDI6ZrSfkR3UzL15R2fr5xGOewyCsC4oYxgw30i6W5hvC4/nqFttFA/rp23OhEmtPlYo89oNchsm
PSfsVWfF7ptSuK9IoMQdkiVeeq1BovsvehMdc2eFZUI0YhOEvS9vUwg3kUgxld/E8YFRyL+LT5NQ
q4MUiiuccBIKu9VWLTIwl+/L6YPBv8VOJfpu0YR7tkLU1JaoIHHj4QbFMbdOkt+qbxCRxlGzOxqe
2zF2RjwlrdEuio+M1dXWPevwGl3DJh/AazjwMemO5B9xTLnSENuTkni6jI1dXnMSKDJPMWUEma4o
ZgYJwiiXexpqDrd/VsW10RmRm+9Tlq4fZEpp3IG5dQ2phMd3qdGVCy38bSt5HAmJLLjQO7Y4zByW
Se/8aYsx1BgLttgVRjj1+cjLcLdBe91h8G3pab2xJNnlAtRc7cVSE6pST9gyWKC/e9462k+rxg9o
uN+b4d/Dnguz8eP9rufJHQkmCBRvuZEa9DCqp30yrqMqChxS5Im8CXyortaK8Pim7QrxNPIXxCyi
K5A4KEIF6qbiq3tLgEU0iNinU1wLeUBc0soEhuJV7XmyPF3JayZMp5ocs+eHF1NpR11lFoDZDJXm
j+CYSvx0oi625RVOsuUNUuS/pmZqYDS1N+Rj494iryH/hYpdMMhftyahYnM7ifT0UP8HJsF/yIdB
dct16l+6umPiGyDiLvP2iKuInI5SBzyKf2Ib7nUdaF+vZz5OSM0fMowwDMKiOwtiJzMV7/xwmaRN
IauJwSSpKcaUvCx9i1JmSvRJhNhXZmkI4QD/pdUcGVhWA7umuf6R1oilG5gMruTeHaRjzPv/VbJs
Bj8qNeclQtdkgWryvfq6tkLavA4yu8m0+DC8Iu550FmOyWPmvlgEBTQCF8qmxsB1ohc8kr8OEdmf
zg4pDmOWPVqS51DoipQT/BnlriCG+z/IlR1FcH86Fhozu8OFjqKxlYbex+qL1XtCTJ77RpMy/QeJ
uyATjQLEO0W5JYnmUKE2iGCGrD0hA4CjqU+Y2DbTxz0pokvn7KPsGGebdFDhxcwM18sve2DFqUIK
KWyUCOVcQ7MKXgW2Gkiuw4HejCMGF6RFsi5ylBniDUgUFCn0byDhVoHB54JOFXK2ZZg4at+kBOTo
9b97Y5Z8DVxiXv32dNgXVFrEbbMN9fue7bIp21faXzFLOMbz1pALP4nrKGrIdLJjnRlzCRnho4Wi
AXl+Sgv0ZEAyXY3Cr4o+WzYuUAybtMaHwRQnTh1vsRp3paelGJ5XYZSVkzX44Z4E1Fj1cmn2rbfh
rJvwaYtSwkkqoLlk/qCubDa3VIKmcCELeSS+oFk2zXZDpoqc78+aJb6n+FDCoxz7kefzmVsQQ0Sq
qlnKzgRLS30M8eqTUdr+LrQyCebWWcANIaqb5fJw8YzUmP+RcB7GP5Mtnl1qpMSELMp+OouzAtHM
0dF0ioilp7gomMKF4ebI1E8nV5dIivEb4NFayi03kgObSHYdBTBAG8uTyHErLHEGA4FRBMPf8pp/
y7du4H+ZSVBEQ5gXfg88n0GaA1Y1r1NQAR4YYTJG03f4qABqQDmEWIaoA3DoKVpjj63NP/tQnxOz
+K2MLy84b1qCd4oON+adG6+tbqVeDkowSYPFF2pfxTHHGwxmbjH7ybgn1KdLOmjuRgwb/XDRO7sM
vL/67cjTG/5R90J90p8yAi9eUhOvbsnxhsnRH2jkmjJy77s24aU1hDxBl9TpN5/gc/u7mQsKfdI/
f0WYHGKwQrtD8zceW0aTXtL3uVnuyL2vcpw2ZLXmh78qAo7kIM/IDqpJU7NFDd9Efkq3/TXcJetF
FeELwx0dWiTWlTd11tAJZVH5kyH/AuXI1PLrt6no3x9Y/ewDwFDZD8TdZbOS7bMn/Mnz1lk0rcyG
O7935DJhUY5/razEK46F4o9SPl0XeJUtfa7BiohkIvhTSbhTH1S8QpLchVzBFRZw7KYPnV3ohhko
njLZiGdx2c4ItNs744XczC3g4aSyI8rWoUbP2TF50ZyQX0P1z+52AZ2JWj5hoP/0LcGFvjwwMvA9
sPqVe24MqwXZ3of3EjbvxPMaUj7K+psn9U9iudvFdFWLLjYUx+gAeh1srCUR7DCeObvB6jLbFjCY
vtULlfc/jjw/DNKmr7FEENOVYUfsKqg7KDniDPnyweZ3/6n+etGGlaPPPdTsVnNOKIndxK0c30Iz
eKe+3QH+onmbGbS2p+CgVJVHDFdkdGdLKN5630pEre8HcXHsnhnR3kjkY3JLzAt+1x6mWNu5DkMg
oEbO4O2aRrUyjfivSzM9E/0HLRTuWg10m6CVI0vuq9gCFf+OJo1wDFm9D6USmR/L0op/rCLjeQi/
WCfx4uOCpucmQ8L43xmVArHgkS31r9U3KhMSv6OjddPFoJhyZIy9d58uIttn/w+jbMYZjQSlocyc
n5TQ6xeQW7GHNZMMJ+qKAIxu/HuDCGOspbx2Fddn0lnG2FEGTh98lQnwdriYZi0BOWnnymQcpgbj
VL9zw8UQwiMCb2wpQ9RiJsKffHYW8pBPsv2Cag/SE5oZZw4nLV7bB1zXXhOejSzzo12UEjSAG4Es
dZAV+LBQcmFjkhbADGVj+RXOAfl1Vi1ZuW8L/CK50pSIAPR5dmP7CP8w9KpUDFmXDmfS3PutK+SN
UbBbeGcUSp8u+XEbKFC8DvdTi2WI4VnDe9sn3UZCxA0xfqBW8ji/ERCSV2bWTuHPDv0QYhyPKjCs
nBsueQ/IvhTHl2y0Fs7VTe2u/P4U4NXNGYUcLyHga7+PL8N884CleqqOmyzw+XYoUiDwklITPXhw
E0RE7VioHgLIJ5V80TF3VZxLu3ey5MEbdLXJxDRH121IIWP00nT4BIOarqyUOAUeoTWs6fzKWKn0
/8ZrjVtc8TpFKDk94KPwiu8D4QwbqKfG4+0RdvcfE6U8Ztf99B1YjyXgakga+7yc7L3Jbr4vz8a1
mLH/C1Gj9xXd/O2fwOX9mpuMgC+awQ8MSyY4AASpuNkawICgkz8dcTolQRVMG4GCuVZmg7Ssm3rc
oOCm8YcZ7CTlbtdSJJfsTq6k1r21pte2QLRxHfz2JFAiuu3wXIdXiREeEbkptDShtLDIWEXXmTzd
XrYNIEtr0qYQfaE4dn9BfUcKSAEZ5HrR8Pkqtsr0+3eikPf1PFAcZyLVMSPon6pH2JkVQLfCTkAc
2tL14kvFzLL6Y0IcebvQHY+oKFmonTP1YtyNRwDYpaLtU8R0WpMXUl+KG0HppkCRoWvODp2pZatX
sixlw2XTwQHgoFxCERZU+CTQM8iV5KRytjyIkX44N3MzTo2/HwjH8afXQyn1mcUPrF+IZPVQ0E0H
lp2FhzsArSufdRJUuh1P+2xck1OAadraqb4M9B6mrb+qMxMo4D85W76rxBjIIc+peRkM4NRsO8QK
0/+jUV9486NInBiA95mz3yV0Mx5yePywwdDUQPxZ1j3nzSsrS1wg9g3RXbIktJ29ysF/CMSyt7co
yHk4zAb8A232t0c6xQ/KShWiyRTNPpIWqgZIo+n2c5N8THe5uPurcW916cjfWJkL8iUu9ESGl3kF
MAGpEKg+60PPiLKuCccZMEb8mhdhSGmafB5SDeVAouFMVj45fE1vDOr9iPVWTAM7JLM2SI4ZENls
qMq9PP2NYoMg4TRgTu2/txMk5SKz8g+a0y4WYAwiq6Gj1UG1pD/hOOsug+Evyov2pdyIVsIwVGru
vzXvYFg2am6hyjCusxOeVnaFQJlk7YaOivLAWntaN7Fdw2OTirookVhASk5S5Mtpcx8iCrB8bBqk
i508LczvkdBaWp4j1Pp+hQRPIidaNS2/1wdTxDfFkpSmKxrKoMh2EAfP4NbNdLags2eb2/RiUVDU
V5i6zn/YxpmEJa7MZbh/4V7ucIWHaCkkkLI5/4RM3Nsi8z+CujQYn/Hv520JCHRuVTCKqivgJFjp
DT1HCUZo36ZskUGbEGZw1pvVQkSCFom0COYWmE9avt8OT+KjXmL9D4IJ+6Cb6ZPhoN6f8ogO9+Jy
OJOeBCQbwn7gfQpgbB4zkEawN3lcbakc0CCx4NSF/SZS2VAjkRWzrhTtB9471sejqsV4HwcxeoRP
4LP92YS9sBUb5zo2zMklY6PdkCjOFCjR+iXD3zhmTINRjYOelEGQ6iAZZINLXVmNo9F/ruKBM8Ip
FaKr5dUuhmIqVwu87QA818Waeoc/z8kEs5vasAy0f0+Z2vGCAQLMPsS/EbGLodXc47baXcOfTPcD
nqOyX4XyF2USV46rdeAHlQoPU2iVxX2OAAxGvqrdJsLEB2oa0UuZuMXbGy1GqBAh107YprbnOCGp
BiCixmA1Q+7AZWVADZH9FTiUsgMjEiifGwDFGPP+eMKVjNBQI4+LEHLGbuWAUYkNSK7njKvKxuyH
qo7QL6HynfmPxS9QsptHfUNO7SOyyC+H3M8GUliIkXT5MU0rmmmvkhV/j+gpXg7a+Q+R5J9vqyFp
mZ9b9tvgXvQM1AFCnC7hC8zCNLEjeRglasHEg/h6WWWx0K6AJyuptpEAPc/KJYc6H7zSGMR9D6PE
jiE6rU04OR/mhRhT9aUfKvjDbx3OLX74KG5+5uyQl+YwMR50yv3OgbL6hNyFbblOhZNUc7+ZouR1
BLajUJ3rLpbcqI442MlY22u8tBZIlpybbQgDVkqx0OUP8MiS1B1CLfCDjM9RR1QmS0oC3YfzTYbQ
+w+qsBJCduME+tKfJcPZhZQmfwATrlNO/bu6LNaycxh4b/dx/eE40J0jvNB6mDMMJYMD+MS8Qpvg
p1zI8ok2bDy0hcEEBOYOYws1EYIRwqj4fsmFyAOnHKZX5I//KK0D6jBfvM+yqygNtDnEU4ARy/9f
4VoVFkpTD/uKKEjUt41f5Dpa1lVNe7xL/yAZLg4gL/N3ZinlNsFE0W6KrrmcrxljuBHyienkAgx7
nUinKPgIprbrzqDl6oGvVZkTEPfQyG4J2TarZtVz0d2p2OzFHgzMRsgHuQDxtaxtaQ4oNZaatJIu
U7L0iS1Fc7zUvBA4rl9Q3e8UDFEkjGvXbyRQnEsRxtJMxG5op3n9U/JilEnevI6dw1/KA/5aL8fP
iIkeo1Hjh+lOm5Xsa5t/1zSf2ok4NdY4sXmW3OI1ApviKhUFsZ9twq1ciYKRGEvCDuuyY5kZXHtj
qaq1Hhe760/s5ujdJMlAw0NTNHFM7jYKAZ+M6y/hgTKKIBsuVZkYOy/ZY0vxyVUYZV6ECglCTH4s
hks3dhcmi5nTdHyjGTzVZ0EoVT0iLWGvSogQe0DMvmh0a+NYVro+C7G32Tmk7eS5+wbmXYuDiCDD
LX8IneUH7FPc89voWYb91UMw00IsFFyiU/taz7DghDJP2+FSnZm0BbMadDxhO2N6DYhfNmdL2aEB
lHmL/Qsa75X0lKbBAXxLCuSKWTXk5OkFwzAS+KxWhfzFOqIEGMdHrypqJ/JuY88PqjImXyu5Zjr0
xIEBTw/toR+ZgeRuhE1ThH9X1jVpQwaBLcQbPjU+3m2CrHCmYvvbzYxilQl1u7FC21/GPgIdpiEY
hQqa5QtVRoT7CWihkKdqBcbGgXpQwoXMQKYrmx7YUrFSfU64RDVqMOfUSoGzdsdydHLpsf4Iob2G
wtzuVbaQz2+TUHJJQnXzEXEwkrzy4x4poWx5cMy3jo8TuK08qPk5YZaK2VTgv8KwgWZ1DeYkH+MX
1YrWLrjR1lgpnWzUXMPP3uZNe+WBStDpA1dybVEk4Xwi1q1tQ3ruHOPTOTeup88q3hCpdvQtowBm
n2Op4QIqUg7a1SAv8g6ai5nr9dQl7S9lKQhezH6tmoZHTE9riMr4enEYRE3aiebLH4IRtkfSCPOs
n5iBJWB3B43OWK3SttoyeS9dNecv2lQxBqndoAzQtUhRhtw3JUrubmV/Gtyo3cpwaHyrQ6sQrj68
bxp4k3d6bseCjp85ccmMGfWOKd9U5jXwLvQDdd4MzjsovVoLXWZWNThXSQnMhO9cJZph8lUIHNlj
tkaVnsgSoS+mR9QcAdwoOwe0Z6DfTqLrW1pH7Qpz3B/vIdzWGA6QqW3Sqf3KCIM2Jzgh09a0M7t9
l7Oql0850nOYyqhU0CJWJxWTCN6M5tlul3RP/JzEMIGcxehyZvpCdJi11oLKetie2cd7wakAIrvI
LdqXESW6eFxqfkq5ev9IbfM6einrLCI9yo0B4DRixPqM4i1exInBQqqsu3/rEbavmeJKCe42SfGo
Ykbonar27PBHY/B+R37nSAp7otAPFnGGXrxeRtbJAzkMDflpQ7l1v2zE/tFMOUbQxfnv2xMMyRXs
3N9n9IqRzhOjQ5bbTu95V47v5QrZKrxZjAR1jcy1oZ8yJb4kRnDeroFYrzYMRtJ88gnV11HDERCk
6XHhg1xiFgbmcf2FyAWHMpIk8HQvPF/gRZaTsjGKA8u/R383PO4JG9qm137gq2wntbSF9xJhdDy/
TiXwIzLt8Ezk29u5r5xNDZk92JBPFV8KyKeta5n06MzjfHUkjMEogYbV330e6cWphSn+fvOPwaBR
8UjvP1fvVgD1laGx+jRPx/Q8SMN8Wr3C7kSZG5NfLlNQKD+w8qwMxLZeJVY1gHO6UgHBdm+xjU0p
qGB7mrPv7PvUFp/x9DKAwdaWlk6ci8sbkgxMMewYop6eehpyEnlAMVLK2ro1frn9GjrTCYFywwcr
8dCFdrY5vUvpNApUX+JVaPHTJL7/xmwQervo59BPbpqJ38mddT+aQww+oseuR0r4+pQZ5eE5dfrd
s6GQYJJ1SdRs6c/NCOMBgX6RCPzuawr5JRGMng3QBFPy31wk+wtnkc7wTrRZlgzJwPaRbuo4lenl
YRfhegvyb2wXL5DXAvXg+HprbMc1vy0U5qMN/e5wsn50HfkO4Zsg4D2H1VUe3GgDG/8lqscEoEFs
RTqGEedQiAzvv71VpaW01+yxkzW6slH8IB0ftI3Ox5G7CbHRBApZpv6cFTn8RZqsKRpQ5zrx4y++
pThs63Q3m/h4ubNLeW8i9phD4GKB21SiqI8bze8Rea90j39CiSsQSVK2squ2FshykBfTye1P3vyc
pwLlo9mQDL0G1amuwQH+QKKtCcQ9JToauLc6cU7zcCSDxGBbZJLv6BvAvNVjOjl1VvaFu474d8rl
MrryO9z2kC/5I7b4nkjBEbNrdK0h4OxWJEFPpJSa9MeVXzZzLOuiecWdWFotgGm3b6PD1vBjADZE
YUJXVDp3sP+Qdo1VAOBUIe/wUGQIZuOO6vc5T0Mkpk3KpIoWn2LGHeZyM4OLxvUZQWcTq7+s4pfN
IXg0qNuxC2cqpWgfAOYlIW13YmkRjOgIf0BuUhGOv5s6Qk40YNYsoH+tWclQRyWqxk3KAPsMg1LY
aVhkdIaTHish2Q3ifeNKDPEVCHeAb8dunEaDV11j/7VeV1etDOZZgOJoBJmzriEDHhYAsAaIiiJt
fimDk+t1VqONGFry/pO1GEpssqbnNuYDE9mVHySfjNlPqd8Ct5KGY64BrnhVKr/DRHYuVkP4enhp
T5B2OZR27GoqLl/3QXYwaOgbtmACgE+X/Cq4nU4QMjglDlTwgk6pivx94P0PFZJZ2/MZ5yBcjV/d
gMz/suGbCEhn5OYtLDZQe2gsrQhhSbnvMgxeKfaJPlOOzAnJ8dRgOoEb9jCA2W3UVdMtpFp/8ejH
nGJmkU0aBzdwXZ1sWtTR5x7uudJh5ZGdl0XmnZfy9Yf2emsZVHsi9dMZ3hTItl34xF8kk+WZPFhy
i+7v5NYOuCu4IzKcdkCaUkCmx0+Iqh5AzYUQZSQGNsv8j10e8qLk5+cE8Z6CS8Kt5Dw+Zhxu5PuL
whdRQx/3G8eH6pMgZg6QUFlyPQspdXQNDaLx+IRGzb7qc+2JL56F2/DYWsECTK6dBuN0R3/tCJZR
JSilA4jmi4HB8F355EV+gTduKEZcgyp5lDiMVOZtxtKVTZsJxqWqWOFQQ1OckQhqnDU8UulgnS57
9etf1GgHoUKuaXoDigoUTC/B4+hdzFIqpflHs6xNeBck8hCfGKkVNbpUp5KDqC/WKW/hcX0kZc5s
Gg7ZxXRebYIEIW2fVhWggECzAHCmmyXAatMMQU40y9uYrqlRg8Y9mUs8WboPHcAP/KPJJDzXleP5
BVXhHUhuj1iL/D6mmul9JcNqggm/VaVYYRBUSAfZTcFldsQuZVn9Qxfso5TzG1v9Wn2jcEC61c4U
EsnQJpBXmY25HL/RPrB0D6EOFqTc1CvEugzcAALFKifykBsCOZrSD+gZsW8wiVsSfEY46+MKkIrD
sVPzbEndYv1K7/GtrjiDcf1kWvPBeH03S9vB1ROmBU0gu8UHcqwLetkYeU6MH0MffArvJKNlEdg3
pQMY9/x45S+k5Upgz5+VBd72lNR5zkPrW0nPlIkOox00hgUzkXOpfS6AtoyuYhvTDeRzZdV4jTRq
gvM6EC21ney6N3ERq5DvcCutdhgTcyoGknWWukKMfj6+52TUnaDxtQMYxZXvhFR28Bsc2dm7ctqx
GJbHnJFaSqXXE3UDb8FcefJx+s53Zd4VlF6ShEp9zaYzOAEFy8gkkfUCmHTwY2PcwBC7+1QOvpbo
KO0u8i2mktIy92gpK0IxaWpHl7UC93S+VA7HL/sfJSzveP30Ee6M0YM+mm5MykxRn7LzLtAGi4zx
P6GXd/gIkNVp5m7aNtceAsHrl5RQHbvQgJX/NJy7NL98SHVAmFKntl96eUQL4g2QbB40YpK5gZC1
TawpZG4Z00pA4sAtYwl2AQx9EISeET2ct4FoGWQjqo+l9ZKnW7wD2sFHLGbqzjCakJCF8num96ld
beqYDzdv1h0+TgCiARK19Bk3FzO1H4A6XImBshXE+smnpw/hlPNCX5w7SsBFACRQy/top+V46TR/
dj2U01OuxbrbZbLIzBADJWGE02t3pp+q9X65g6PibvrSBK0KT8aUwuUDKv3Z3hYN5kT86QBC0Sgq
bVNEuj6cu5pbS+DA58poconKYp0AHrOvSjqQcWQyaLCZ3oPTEXC/+li+iC9wmGVIkoaOnONfyK2L
HzOa7eoG7mzfCQsp4CF3GueB3yyHYIfGhlRzzLGM1jfgviEZ8cN3tSOLEOcoXeLkFgn56JNtoaCo
rtxigx7wiHfp1aTVU1V10QI8NNhUKaRB2xrRRttyI9TCncxxp4Ex/Xco68YWcNkNI5tZ7exkKp7K
vmDRQWYnSe9sLg8ay2m5prqcEVZHm8K2xp05OmDxYxXJnSBS1B0M6LqZCVw1vd6f2cZmRK9OBBGl
cPv+N2xLfS5eNuJ6BP7AJRzshnwMzEUJJgmvs97s+XuVzfb4YtLy8Ma/KmTvKDHoHgP7B9vJgqWh
AL1c83tfXsyuU/hGGda0PYvMg8uY4V4GXBDNhwSacnflOP794+g5Bybq0TUXQV2ETRY3Ct1kIQJ9
ywC/hAcUxDeyqv58i08ZE1//AHYUBCpEIVyFv0ZK4A0ufU6uyRtAfQFw1aE6WWPBfnCL+Ftv11cK
7gnzH79pQ3ZP6m8RdNBCV2tGrKIclCcpRTGAKOc/cbqGH+M0Mnw8ZglxCWe3N78FOhXjkvOhs9xV
3Z2b2ku1x4oc96cdLy09M0j9Myxuy8PWWkjQgA6WFErPnPj+8n+p+1mn2FgDiJRJkajz4VpBHBN1
nQlPykMu2/qu+GVEGOodA9+mcrosWkbvhalGqxmTmmislrP9WWEPrNLw7VqeFaM5SJsi4ymgaiB1
jhL/ASpsXY8Beu5Ik3C380y4bms4Bori19wevj683HZfkxJHvH6zQ9Z4hMaJHZHz0lXC0Rt5FZcI
XQ9ms+Y7EhGIiToRp63cBHBDb0gJrGBFw+fBKYW0WcMCFVgjKyrR7HfgGWypXj0gsh/81rHaEfew
8kPLvr4sDiZrjyrLgJb9+qLA7wvFPQQC0RoLJ07M3/5BayRR6+9GxwCTRxXTQjQuIng8xCmy/mGD
XOgslCmKYW8S9UjAxd5kquFtyD1BWtRe9dZ4AQAZm0GFik0liWzCEkomR4zpz0EvOgGmqR2Ruix+
P3/5pFajGCLprPf5rHKhyCFXnwWvsi1lElVpbD9KHWqLltLNFSeefTr5tKtku8dlNMUXPA2YyM3q
MflGd6zwEArujJhdCfs8z3I5bwBrU4Kr2GXGVCI4zrXUhQIHEygx10D18YsN1yAVkNq4oubQT4VO
xLSl42iUasB1QrP1teLebvsSAVsohVMo1mTL31Zkd41JpLTtqJ5ZRvrPqEvO5JfZWzr0xPzluC7s
FR2ieGJUUZwA9FkpZ6MzNlYp3juvDnsHkLYolGybAREhHu1rIR2NidDCWWwyYwtRimPVuJiyZTZb
ZOAShBMcltdaKth1rZT+PM+mJHsb9MDT+7YKTK/av6jM1SBxscuJwQtTBPq9EtNVICdjMO8RWpFl
t4aUIcfw5juoLdwIrCbPAQX6flWzOMIvViOeDJ/t4zXUXvBvn75VQWLYx0+VboeyzEWvAU+aWMtM
IvN5Ewuz77SK1wK94kIIT58VqzYTELyRjH2J+N80UpapBN7tMaJlkQ9pY1HfuYXaAM/vfXxCPFSa
lEVdnHcP+g6an5FnsWo2NSf13KmxmNQbFRzrqGXZuXIKipAH88nkxv8w9p8asOT9RnZLsWEyksBR
f6VY/dJRvr80/ePy4TreSKae7jZ5WHLz8T3ZdV779ATciFmZsjcnq1jiXkmFzj+9v3+x++3HaSsW
nm5zLESelDV6YIw3XIxJfGgKuhhuQg/qoJmOUFBNFkt/XN8m7MK+5Y3qGL4FaWT3K4zUPpoP97mi
abKGQZF8Z/g+eNWn4PrYAo91Vn1RFYAKYSmL5+Ijnl+fBuPEwkivtYcVQFCTZynmN1tzVmvfYf0f
QlB6nipfa5tD7jE6Hch4HbKjQ3KrSz/hhxD2YQqxLPY79hva0YvcOa9V2cWeHEa3Q0vEriuPzEfB
VyuDvDnYXtlQlhzTaTye/scAdtpiOc9JsFmBL+9gqeWxwPv3BVHKpZGYKQQ3fSOeKdM0Ni9MC9/k
i0qCrmhf2YdrxoHISeD+pzdzt9fzoJQSLf7bUFDuVM3zCx6pAARmpVybPGKBT1D6YswOKpZ1BaGu
1b1G1iHGhy3FDBi9eJnY0S+5YCALfM2eusZjXi/NDLhLF2ca8/xl/qaUtDDqMVgTx7mocjBXkT2V
fxEjdbyNgke5Dqv88AoLrA37BUg8/SmaNRyz6uxhxNjphZKAeW0d+z13K3Pxics9V25P+kDQXAqh
VwvYOpI3RvJAor5OHzr3WMij1W6QibpH3k0UpjAXP3CN8w8DiA6AHqkIYLpkr9rMXRWJA36rUdz7
bN769Uj1ez2rYq8fWf/2XPND2jSjOzYo5QFVCEDSr5p5QRDKYtULZbgBqjAFa2W2Adu40bxRe5e6
IVQjm3kcBiRra3dSO2sbUY9EyLqMUO8MrfZWTForqip7ZFOk6D1H0ezzoVXeisYdlZ9XEahLzhEy
8B4F2i7TfZUu/xwdLNaji13ehZrF3IHOn0Ihv1bSqvq/FQN6UPjsqvE82abKP8ci3NCB8bjBTK6I
58PWTAHrtojL1K2N4QudCSqjfDbzZb4TcT6fT+WN0buC8Vh/CDUvDlxLifJpGEVa4YYdoO2tptz+
MBTRL8fYs6qxyxNLtWigfi90aifQGnRv+X3KiLuE55uQgZVZeUdQSHmZ5bRiHnxQStMZHwIae1im
AR7LWNbZiyl/JmUtbHNvHkcuj4qRt2XFrRGKFOPOLMa95BLr67qX8RYoqsXGQuSSX0DVoZXuxLjb
//b/+gR38LcbDKXyK8tPcKMYSvRlWKdqjunBQMPCaF755Ju6OqonJWG/aiS9+r97Mg4OZOblGLZU
CkyoGOL/QMM60fe3eccBFwF/IfsKcm+KEbadWxk2iyx9hOCE73vAXMq7aKK8H7lrr7YnwaD1Mrz2
9AqYMRiHHZiNKFyuzTiDNm+OHtaMnIGMdq0Q4AT1jzotxAlOxv5JxSGQOotfc++fZnK3mbnHIYAH
5pEvVExvOJjFdV1JHHsMeQTLuZHvcyu7Mndk/ssbL6La2yCR2H+w6q3L/jHnLwHKBLVM14PHXgig
XYc82DR6e6bm2Cu0FQhV/2J7cZK0xolids5ilACLTG6D1E9aiWBWVKrF5a0LjgwiXnPxv4wK5Yr7
yKHfnd5/3l2d4D0pHXPHcZ+y8QHJdRocKuEDfygFmFqptoWLJlBEf+gHGdtP4vh0YiG2DVS3onH0
JZPwe8oWqj7YEQIJWdJurQF3sA6xepBMTNUsWTgYh5Yp4+gx/PSZlmIPT0570uW9iM2bgPuxf6HL
tefn+H0qqi9fxxrpcNv9JjDxPAwP4L3/WEia9OOxY50i4by0q39bsEQqbpPfbetZl9K9ouww6xtj
3JE+TmFlLrHpO0b9ipqERvp25RtOTZpY0vU1zhlpBgYf58DI5QBo5nUGauNUMMqhELZwUvNQ3Wvk
EyLQVlJPren850qZrZSYUMBl9so/s4hDYWYRGXcRPWCvDPpYt96Ub7dr/seKpx9EahDOoqcr6qxc
RAxgnDaBDAeWVv84LB9ntGCNPpJ1w6zX9B4JmGG9RZaniF0A+S0CpXr3BtdONVHMdMNKvtomZrW0
liWhQ3Lyf11gCLD+YdeT+ybWebhvdyJS2PtrH3oYwFUEbDBZYaspqKKISQ5crl70yshshPyNQ7+A
qh6XEj/8hv5Je9eVGYQF2hyQZI9ENlrcP92GDM9tz1WqcdVOy1dLhbKqia3FGjNKZvl6FDhH2co0
++ADR5Vr+T1LTOA9P9/uJqPrUfEbxcoI9AB5nSOZlc+OMwbeJPfZ3B06luVMqN8rSv/qnwlA9L1J
6ozH3b1UheUcMjoGKtBHqrsmT8Z967Ow9PCzADJRfF3luXvBHhepVNNWAeede5cwaXEmYjHAd4/4
OvwyjcyuoU29VsKbCCagIecg5bFWzq/lZDac6wTmNGlRIlLNYv+gGNdrSazfmKgog1QWorvaNg+f
LlK2dal3ogL++gk57Oxgtf+lfSbUQvHcAgDH++Kb3j01Djk3iEk4d+CIvH/PDsQbhilaY96EZoJh
sTpxD1zprg8p6UBLKnEXH1cF4JSn8hI3+htr3blKNX56GfeARU926oDFCTibbj//+kA+fTB0BfKX
hCRQMqFPQ5AJI6thbZsjAOfD1GlOzgFGhllkAMINIGVCE77U04JvCMfEykmN25SkYcdehTmeDlwn
0/GcY4PESeYufVBsAggKTyS1tvNcSmeHLm1oqhrib4L0id1Ah1GlKoMyLkGQayebvNDeR3JmuyzD
cazUB5DyBzc6VMontOlsnn+/x5ZnrDdcDeRnEqYRnBjMhTlKlTl+qCh5qmsEns8tSVkP3UXJRTB5
lK/32vKhjD/hbB4EF0DEIEqro+T6JwcA4CDxzFk+qjq7WRe+fGIzO/ugqajYO6RnKFRHQFvEUYP2
z7E/8ng158CzKs/opdKtGHOyaoRZyoc+unmmaQpF6r2vAZXnpSZY5YuwGeO+dfhaPOARmtwRWhq3
ejNeJv4AxmDRMJdLPBd6Qt5ZiTJwHgZJ3DGnpwkTU7zxNSNoD1YUE5nK9skDTGXaG5HHDRW3R53o
x4F+WM+uLakoumcYJ1EtzSAbIf5SvXbiNDCAf0HFsAKd8wLltHfuzDHI9ExPYdBlU/WYhB2SQluC
qK/0P/u+N35PDtj4NBkjkKbwXV88E4UDr1QjVYLpFc+8JgkETA6Xe1CyfSw3wGWBgj/XtInkKEpZ
Ec2RNS5UWzwTk8LxjM81JfYweEHkyftNv6ubnPcTFjB1qptJdABimaiDE4DuAbPXp7kFywMNqCn9
PI9h+IJJgcbayYGftB6qZXGbuv6NTvVK8ORF2zV38A1OnKs2ZygxgpSR2ivPW8RH82h5AWBBWhEt
gx8YvWdB3I5y+qGT9eQSmFhQE5jNKIp/J+O7o4CQh47qqlZO/+34fTBomx4QjYfh6qh1iVzMkNOk
9GIE/WNeETcrFn4C67jUMrMvhnaNl7GpQ05/xPSPWdZP+qt0keGX/m77U5QiJ7AsqDD3UIcp/WFs
/KmRzgj8igf3YBrNQxwbzh1ozK4+vjCx25Mocwkd7OVqXaA26duoKSSkPnwm4TH3ZZDxYRJCf12t
j90nWF3b0qQe0wAZFfDvLOOuuGEm8p1yGKthyBqxc9byGWvaI0/arZSgmlURupG4TUzdcME0IFyM
t0I9MfCOPI4crt8v3Vnf8WHlW8vFMLWwdyXTmJF6e0CEScchdf5AbL8/XuIylIOaIjvHN084AUMK
daXkMySdvBvWmumNsmiUYdK9sdmOBzH/7yBxipKQHe/fHatWa5kZlO6v27UnIWmaNOLHH1OtaJwJ
ImYtidYg1OEJm6bLBhEaHVEkfVrYD/FJ8g875djSaNgeoH+IxAYOF+awqbfO90zju687+zVuApt4
ksi2lEAWP4Xrhb1kWx1024Zbba0+OY03Ufyj3xuN/4GkyOKep+Gq7vYLNiT9w3pNBbDHLoZTJQOx
EZGUuY0wKQIZpNHDeJf9QNmdhn3b2HblP5S9q0GnuZ24EtHvQOsS5uGBPh0Z+s3sdGHXJdgSWubC
EmxNCmsBEbuYYGVL4pFWXI/zi7sAlEa5aFDrnOb5VJmUoxC87sp8qmrg9UQ7mzWVPuiv0KF7x0Jo
0OV/LtAiXNuHB4NLdjZuRaXJ+CGpYZwL94YhcR1ULJFORAiWaQaLve4v/6fGrNczuFMjEDPWxkNe
hZcJM2BnGBfu1dl2PcjQKyzG4zZVS3N8uYXU7dJGzgadMF80XTb9bsbz2ahW4CBjtNDhaa3tmz+t
bp/IG+Swtyx7LmFaMt/VpLnYFURL/w4CghRPtQOZc8Nj75y+nV0+TCCOHI41Ygw1EZtXcp+MboHx
9x+lANNQLd7Y1pNILN3OGrENUfMentTlD5NVBpug0dw1mH2m5ik5mLEgoLnrItGDOMQ+NGntjm46
BXjYzVRk3dhZ1yUF5JHDGgEiM1B2CzENEZO5aVOzn+nadgx/txRrm748/INLkQ+JQUadJpY3I2Ez
XtuKR61IRDaUg2ytBlF1hsW5D24JlzQqwkKK3uAIJR6enLyLBw2Z18f1SLWccdUjCGFrIu/811Wv
a6/CALZiL0kcKoYnAy0UVOiBkpi7nn0uB2HCcV65PdDIhosLUnoh8lP/ZpM+8jOx8QUmX/olPOSx
x1U7J3toqqVNSDHftOIUwPIZD2YGst1D+/O5/0A3spAHSaEZzPnZyVVlKWY3RKbXRcA8pfq32IGo
I4RylxO1cCjrd31iFx4lZ/Q3iRMjzHLMr8/4blq0+u2MliR0EVJJEL2ZmTb15Ke24TPrs5J37bNU
RVmQZ7WvaIQpOiQ1NuQzoboULCfrCPgUpumYzeDXbWdtc45bl35YBnW2V8+MeOCGaY1XaVqew1Rn
a7sUuqYaXM7XBsdTPFHTV66ja6xr/hK240zJlCApn2WRbh19HD3ylmCrr8UQzM27etaAVBQQgsYX
/5/m5ZpJ4ncHTCOfVDop8ZF9Tawd/+4OnAora2zMh6MajpBqlOHsiGpjUdqYPXoquQVDiCU85XJK
dg+KFLiH64T92tp89yZb6BIlL6TtKhx7sJ2v5pmcZzXOAh33b3D1AurDfHvYMNZPK4I94qSBIaJd
gjckVhMCHLzkAmF3Y6aGuB3868pzKRF05lNY7xP+/k2/++3tBU104eYHzHsXxY8UBR82c8LMQ4p4
PGOY0Ydb1WaGpAIkwrrV+JUGOt1HrP3qElclk9cvhwvwvEYiv9+7kEqLrYJ4EBJhHCqd2USjf3tL
fe6GB2h/fLNMCz45Uxt9cthzJ+F6dBzoS2SRSP91wCau8PASXCwM487Wg6xlVIRmaUhIpholtX1C
1I9d+uIzbhUMHTo48rHWT4jcad9nsFVy3lnFlcsp8E2hTNMRUggg6mMTGjVmaogOCbvaOx9jnT7i
peo+ojmwzQQvuCn1mh0F1mGEB0jeUYftVzu9+musJVpZIxQwlvcQ/1JO+Wo1GvHlNp7dAxCLM1Yq
mxYaYqpn/9Huv+leeQTLDJ/qiq6l9SPQEF9gr5MTa16VTCHq23Y0+1Ai70dPpUYtIS6LiX1/qbMk
jk+cLOwgupd0jCcKVPhTXZxXqVzz92bu7Th2RwQe/mTly8zN9hiA0Lkr1CX6g+5cr7sVr1Wpm2o5
m0X+PcqiQQpWjBKtOsVL3m+xzsWU/QVrlr6oONYdyo16rL/tDZl0AxCYha6ZXkS2FoQ+UIQS9ipx
9VtLXKCj/vxWo9157N20OtNe/Gv6oEVUWBRYIYwiZ6EoqrgztsJgHTsgBp8+uKIsIaU/8M0U84g6
qtWkLaBptMi7rJAc0jYEsGvGBMmuUm9Hdqeamro+V/pGLUGpiWnykaGyBQ+zAUcLZPqKp2oXlOWT
pfgZ+uGjJKw0fJ/5mwYu+5gXI4LN4LvKagZ0kwF2azElZg7u+rIqN8vTOKUX3d4JiJLmyPsYLJbU
S0+LHcqElheCLupHZVmyHUiNlU2X5hJuXuEdk4XqkDGiBlxvhDvWU0BoGiwCDTHSoQD69iubF5AE
PnZZz8LCyyyBG2vPhiqJmZWkX7xOPEfwZAqKsFah6e5uiDEFB/JiRo6JeBNlcRjpv0Ke3sXB3KgZ
8OknPSnYfeOMCetDq9CGy3o72nkQhVu1EXuGZv299ldYhtwMsHrB/Uf+hd94/LLZPVxyYDdq0iB3
gmcHhyya1eR7ixDqFjQlbq4oJnWWejbUQSwc3NZHCLI12WGpqS7LpMqvCvZ6n38le0LHvf1AV2IE
lzqgwHpKz4GT2q0rmS5QXLjeLRV0LNNcFpQUYKA5DBEEiBMwJVsKBMo07DdoG+6K8uF7QFBXAfSM
LgWw07g0Sg6Eku5ngbN8Y9wfvqeb4K2fB1+Z5LDiCFjrrqf86ZK8zNtf/K7siCB3FgPLWdECfmM3
d9nPfueBa0mUEBC/MPToW7OpICU0BVIxUOqYg3MqIuRrBRHXFLJgszYn4mlWaFyUyLxsG3R8cb9R
spgNdIOVML9vuRYgW2ctu6lXOdRs1jVVengMFysIF+Whe4uXX2GKkzxtDhP6KETKGsDckvMf28X3
ZkVw8+N+opxsJJ5jeLEGQDCstoNWfQxmESWcE+diASkW41iKpgnTX2Wl8/7ApltqwisFC+/V7y3T
0J1/CHiU8t2DSV1fKWU73Y5zmwoCtzz2smkm5wqugLcm+uJuZGB25u1m/aSO/r9yn/vMauOTQujC
9ZTRJzoPQ4dxesndcbVqdhgJuh8INgJhiHGSyVA4+72QFk3RaLjHuPndzIowOEdtV5Br/aqJJioz
quy6kA+RaAKAeFa7NkkzquP3MLiwEEngi0kvuThrC7NAgVlcrzEB8PTEw0T/5F8DmgbiFuys6SML
98ffzZZN9lYN8uxjD6Mz+Gp62NjJxMurp+FFhLsEKnxTvimbcDukgLf8PcYEMDJfElUFnf0WJ9O9
TPsKokdlEwaBRpm/oqr5MiDJkQUtb8hdxV0J0+zQ/e4CrhgnrJkWgj/JE/HQt46HSfStiWga5Hib
2KLPiCT8VGM6Bt31Y1/JLxgy1EKe7R6woVqPFTdA5q9DOAZEAg/GXo9nFU43h+7uYguu8LxHxKzj
bUNxlfWRbFVVOTrZZSLxgnuGcu4OLD23Sj5v8hNoM39wxx3kOlHnMXDq2f8Pizi/Az7PVp4DPu8W
1m/NJWCrUqSuIKv60gYsQO035961/WVZslff7DRWsM72rWtmRaLYbIFqA1i1JhEuPDj0FzSkovyF
Id8yOz+taiUxWkrX1u5IRZnoSQKUvYsv0+CMnfCOyaKd2XnhpH1sTL3bhSS3WWnKeiXEY3gY7aVA
o3kS6EPIyNL1jQjn4lvb86UxNlRa15zUZWUKLZEeO1pBahUMGyCVcqtz4pYf5kxBHlpTuyZTl7rd
Wb97Zab/0jE0BJx2LhIRiCVMvKffOR2wI42EGVgNbrJweWNcTFKcEtVR7kWIqQfAiiqZh2/LCcXB
zt9TydqVcTYnshWq3Dp3tH8pjyvojEkBfYQt9qo5j10hLWmFrAj6HNppyYo4tE+qYWB3tgvfqe5B
O+hJOClztzgxdkRXNpavgafTdIK93nke/Y5rZwdBMBPE4pxmlk+SuPRjScZBzrhE8iDh2ZAx331E
zdJ40kEww0bFSYWspgzwxdfq0D0w+rf3Sa6O2Mup0F2iQ3ZzMdbj6ogSKfFCPbdUf1cS+IlHHcDQ
xYdso1F5vYZxrO0b3nkFIDcySbCZICr1slFaXCfI70fPKUyPoxSZFSUn5FgAIyxDKllgcXP7SwOY
aDU9YPWaMyscfh2+SiobtBtavi19xgxiz0FGdHXZtN+z9osxPhMyAfOvNY5fSmnzCMDqw4n5K8c7
7Gdt4N/7E2+tN4VIKNl6MxGQE23j/EFcqgyE2ewg5Gp4HoWYw78Ue02DiWW5QWlE56re72dlTrKR
Wo/UJZwD37+Qv9OafYu9HEb0u/YLnVZNokD8SqAQLEWvNUzsfy/SPtuZEy/MFUbn80pJlFr4zet/
zbfRsk3ElzbiD2CeCRGDGiUg0eu/S29y0PLfYIzc4FcfVTAOV3X3+4cJ3C/ll9McvDF72f/ePKRG
bKmv+/cC8/ebZBBGTGFNm+1VbliYZq0JMepC7rzohcUJM/2HSi9RifqrX310w1ttvMjRsl7k2BkS
tjhu7Ms0UjHptb0e/MAhxMKrzuS/xuzEjJnac8KUQsEb6rIdk3dVG/lbuVPTpfDM0WNsPhc8sYxQ
rPH/JhnX0i1ERoCFKZwZfVmPQ3WlqgYgI1+ht55P3okAs6+SzR9KE9f7p4FgPD061l67pZHaMKgI
R1n1HOL1U9KYu2ThH1gTP/ATaYEWhRadJjRxam06sUU3x6b/Evgvru12elQp7XF4d8A6qQOLosCm
Rbv24QO+WFcKY30jVVHBvMtUkNicXk56v6A8sYujz+zK3lZwi9ZKGuIj9JbflBlSqqpQHJXcN6bE
99+yATRtT7C4cbVy+LlXxoohLS6hQOqJRN4ixQhP7kREjbhKwk+N1AjrT1kE7G3epi9rOrRNjeL0
bBJokfNwdeI6mH5Vfh1XNJyF+4S1ATl+35jFCP9lRdKAG+2F/X7Z1a3DMiJhZoOY1i5wrZUIxdQy
5FTkVAhJqxOKMxmYTHBPAi8r51mV6rrLErrm3+AJ7JlB5CuLyGUwSxT8mz+id1133m5+r+31dMM1
9dsM1YOfKZjgLwVcZ7IEq/uKSWkfpocRxInsrs94mziMrtiduoL8q2G5VYJvYHz9sYbZrp8tl+UQ
KGdAYs4+kHco5/dwUO1CMAltF7JGRwT+XSEqaroVIrUeVqiIRnKaiE0pZ8zbTusJTQWdmNUdmLgp
/KlMLd758o/RAD45msClX9ZLAtwxKNNz8mTSk3RlzbGi2bL2cQTGlXkTIRYlQHe84HBhj0z5ihjC
ZYnfpGhKpxs6Pt41ADXU9ZBKu/qidW/ys4o4/1sXXZeDgFjg2ymw7I6wn5rSmTbYQ4y1Iz2D0DYa
Lz9KAV/euKssI3lAPbM1HL7RIGPvOVEPfopPD9Stbjs2RDLu0akinCy+dVGPsST2l82kpA6T2fhR
lWF8nW7qNAJIBSl986EnEvEuAC6DuSUULnT+ByYInOGUods6eFXi5YWcC507PVJE1zI4luoKtZio
Jqju8BZMOhNYGSqBTcUhcF6BI+CTaNA4CukFx0ajC3y8Pfd22mHiRp2cR2CkUDkdmj8iqp2ryASW
1CafgEBDDHDiPA8HffN0VnhBpPo84B1iNYW1zUQgcTEA/Y3HruW+WXk5bkglqDwDWKEuykwJsmj6
zGOaimLCQ25I5q1iDKCYlcBkTHw7jGOwn8vp5dyrYdnyftO7VKbVrcQoeNrKkVAGtWj+BrsaudnY
37lzmZ1efaBJdPL0xSRRfdW8kedBR3ObgXf6KAOOKnSgfh+ETFCpieoqn8jzwoTqm0tH3B6KH3Th
1qnBO0vrIP+/lwv62eohEEejgVPwUk/KSaYVgBTJnUx5FDXA9VSQABtUDxPgyE17DJPBxVCcB4fT
o2Cc3AS2hUS2AMBdK5biIMGDgkkRUoWZZF6sF+p9DhGvWrw/sRkWBtgHM8uB21DVoqaS2KB7SqTi
N2SO2zX3FAsUFQkdt3mv7oEv2PWfEr3MVQlIGwCiATcyJc1a6ML0e+jSu+C+Qw37kwT7EkbKOl0M
Fs4BO8oVMLUP1jHdpsnQKNjmMsrF4JhNjDHLk8FXrG+vFxVtjHM6JIo4hZ00ePGNfuYV6C7lM0Bc
GoVGYQ2a9rn00Ybqhtu7DRmhtTqafY4MBOKU1hYyn9ZdUphCjlqckzSJllgztajShab7L27Uw/Jz
CbNBQJGHhMUvP6jODkUfDGc7tS7rOD/o70wIT49eWbEaPE841YcFR32KjhycbiRtbo8543pvUuCU
82/EgIuv6X9WrxZn+4fEkfOP5rLNNunBvaSWXNeidSQKLj2q1ltnOa6YExvFA8O6YigwlGcHBMek
HcFDMEQSD+aKTvnlAs7tnhw/WzDxm3yKi+lD1ZEgBYh3k7RXe0K792QuEgBaqA7ency1nklQdanD
783kmSyCcWotlBnNObjz8IXvji/ny9SO/OeqsHZJgbvyhbq070UJxC3GYy6lx7Qmqu+BcdvR8mNr
Ib9WWIQgss5LY12S9txfyanqqLY9efKYVl2JDbIDIoOx+7onBuf6dHqyQQ6XVXuj6hZJc5Kep79y
/OXa853uZoKw0aElrG/ETP0PhdbvaZkkFCWHcTSHSV52H6/QbNvpOd73fgN2mDkN72JN8BAe9hk/
6BCd3oGamJi2TIAMsmzF1LzY3JJrVtgp3H3gtlK/mBu7STuxqb0A9UqQpM1E5/gfMnebnrxWZpKY
xDw400+fXjdQBKLgQhGAmJiE5qXR9kw05+ZGrcKoW5UTOLSpRTMZHlSqz9xzndGa5zggOt1FjavE
xzjKY3qc7wreovLPHcrxoqXSVfeKPF6R0ZF+wAR2JM0rPiZxDoUar+JuoMitxf2LWY+llZMeh2m5
KZZUqoLASlO3f9HL+otYPIWbevQUTw/S5bj/ABdg0460Nts7sucsCF24VsiLOIgo0jCAOCRqDArR
ow3ydZIgOkhpfKiOq38ER8azuSgAaH59UqYLVySED1kvSrTK3fYvlxXMY5I02dB29BiydfBgtWhw
/Jjycvk/A9e1hPpK8IeX1RRJg0rzVJ+N+5q2fUmavBu36givMObP/ZlucH3TesuSh38JNDt9OuBg
WuQ6HQX/IhlnFgFm+RzsYLVQGCBQ3l9FuReq1cyWKwihmpGTuqo6s/42Q1EcA2y9/lKaZLCfSlP9
rfaLtgZ5nlPeq5dNHtv80Cysp4QrpjjLCeuedjVfJb96ZmI2ZgoKMCZGFMghztHVxZF/JLgu1pWr
QxNiRVOnYzXYaGMLNwxRDkxvOVhgBExGbOXWof0m55503KsZlu9CYRm5R6YrFrW1dH7kIYPfQv67
wIV1sriYJkxYb5AEpDu9NIBKU+Da6eSyQbcV41a1zljUnNXI0pwnFH8e8nC4SrIXCtCL+DUHFzv9
CsBu9icF43El90F5DZ4HAxeIzli8lm0NmyXWuRFz8kWQkQMbO2F/GnQwH5TrEK/k95mqrDTGZ2va
1PLYBlQyMN1H+0Tz27q3d8r7+BHzaZ/yIdcyH/G8VzB2XxpPtglht9u6AN7jAk3hnrboTBBBMMC5
VB8T9GSQXDS7mTzh6MsgOoFYCRel3pDGqBji8aiZqVB/F6ofjhzNPxnkOSMDjpEXdJx+ORnnjRto
uEpgmUQX//rzcz/587NYunH5tUo3ekYBCFkIEpGnGT/RujMxgW8DH+qUaaT5SU7VjVtvIbAmZJ7f
+q94hTdZSq+W76eH0vlXNDBomwBXfmnHyPY/dWqTZfShF1TX0e4GGe5hjF1krG0K/1oUhOMlzEr0
UsMz9dGcwhv+6FXdWVTvsdT0cxgBEUT2Ggxe4sxTMRBbVEoT4ZHCJYHzQ1BJdEJ1iHWCGKGKXE6A
iNFdz5MCr+n/aUUKTf9pdlNV6+yQiJra8teFWfzWRdnX2W4phN02tlD/L/3otDbFW6fxq2zp9XCl
kabHk7eZ5xkl2JN7+CVEki83aBHijr1yCBg1dR66J8VhuGSH+Ew537hUpEIVg7/PAjbDgm5kT+gW
FcVN75wgMRVnqB8KCQsXFqcXiYPCnJuvUekWaK8uxxYFtK6xnsHVwUgb+H4yU9CgUCTGLFtgCCsa
TevGy1IUGjXgZM9DPdLb6abAOVUKuX/yjY4OU8WpmsQpmnHGns/c8j/ryQAtcXz60mpmTn+EpUHA
zEaMCoOAz0sUcpk6jpybE3E6W7DE6n/0bJ1QLDgYklkmdWadFYdsbo3fw43L3QpYiHeFwwNfmG7F
ocaXutwpG4bofIRmh/aHBycFyGXtjO99vBwb/MhwSXKZYrJsXxh19FLUjUJGRQFCcHrZPrIf84lX
zmzkgTbbIJXOlQLpAAfUM+4vKJuCqDf+/FUOx3rPPYCpPiyvaotAZ7lzzOJGC7sv9mP2BKn1sHcz
KiQ2WOt1Mbbexa422I7edVDTnXZNbTf7akgM5GUAomJVmGsMPRRLKSC8CNGcX/culRTvfTLjf6Pl
DDadtJliesnBqi5E6V62Q/rVkbFo1OYI1lXeswrswNm91BcYHgzdWinWdxNTISDgpy3F4hq6878C
4MVjg06svwT12V7PwvDICgwZ+K5LkAE/NEl53ThFntozZQ88Si93KPy3QRiJLLDp8GImbBbOL4CS
qOVDHVMqSdi8RuePMuv651Nay2WywiZj9p+bPj4FU5482bCanUAsbIuxNx/vDFOFOTNd3lXZParq
B2iYDHPxYWp1AxymOB1oYtZvV4zr/GOj7joONFJT+glhj2c2UQ8MLMUZVsvtD+PkPrFmd191YsNg
mYsVCEvmAPveM3Vklk/jpeCSg8qViv9UsolzTdDzHHRfiKgcMUfOTRJnka+O5JjwWtpWJw8WKGe/
J/ZXPkT71Tk2x9j4Qft/b7xP3tUwe02WGIFfBi18fuBDh07RheNrzlwTr2FH8ldtpHvGsjjqsPTs
sTjKMN+ug7hX7XAbEHJppBjc3V9SsC25aDL6B37YsUS+fPHAWoqsQDdYwx6n6Ksz3mtzzG2AIGQT
GGh9ORqoyHIeBEFGVn1ZVauP0osBd2gki6m5BbT0xarH5ZUQVZHz23rRvk2XPrzbaBgZdWKqnjrK
NXmeFi93D7jpIrt6xLW14UYmdYA1VwXDP9zI7hJG8RCdKmhZ/DMG/DMZALSZpL0tCn2QY5v65Mzu
8KSalYND5RUZrSoDEQfP7IEuZ93yWbfEs8+Z9GgaV/aDm0zxn+gvB5a3PB4TuQu97vnrFJp2PTs2
U8k6W4UttFUXX9g57KrUe1yXEmTIUvgMgg7vX5cj4+483C3UTtMprpCm60eGO3wYKrI2Y9BuQhzV
3y/xuvurAlX5QFNAbCWoi8nOAHOPlpl4J4xaeVbQK4HTlLXybtQrw9FWaguKX2QAWVS8SB2uyF9+
zb4CSvBfnzssSoA7J4oQmiSE1sc9LY4t4wvkiIOLLJ4FUviVBv7cD+/pjDJ4yWltbbNN2kUgQ5CD
YPUZPjSILv52hG9JNmxS3o+lFD3dT6bvISXEn6vd7pVcO2b0KECFoCoDGaw63jKjBmbwFoCmPgk6
+3BUnNa3r2sP8vHouMfsubdAWU7kh4cdMZjo/YfXfzH/UdyVYAOGOrg8/Wq780RAOSY0jzIBi/Zs
f8FUQgsPowiobvX1jtWtEh0IKx2boWR5y5gQQatb2OQCz0lqegd/FMvYy+GYdrxA9RttTC2ibFZv
Srx0LWhvzpqHxo7NjG0iMG0szzEaerDdWMd8FO9JKAGMJrbXd4DmznJnPBzv8ch9Os9Kg4TC9e35
sA5W1kM8/P5E2cPOt8Ixar3eFDLT5VKWWTDw571RDoDndg7AWjDVwUxjvmIVpDB2eGuaxMoZaWil
yG1/nQ91/CXy2kpKyRtwN98jE7IgmUTJ7SgFu77JpFCaQQ5NbvXIOrqa4yqYnP4dF9FwJi/FtbON
Wk3B7uLqcHqmsEVPr0qchC8TA3uDT4snL39KCNQaTm4835nuteTkEVAoJoy2VtXO2cgkFg+eftD3
0qw7Xk/VB57uLGgSsKGLQbskHpvMPnkoq0UamBf8gH52YMU0zEgZY3JuovnFT8POY23uory9Xs56
rzLDU4VY/9H3UNsSgC4pMHchU6eR+CgHoaK1AWZlHYJ0XmXKzb0fuwBO/FLKEEt8u/oR5QvOwHK4
/Z1WMcfkPHAI5fiX9KV7jSSnvVp6sitAZZ4P6ZuQTfEAEyqOk0adFF2PO6BanMEsUkGRSDDpEvzX
d+S+BFfiSs5Fw+rtFqy36yXYw0dG8AZ8QAS/9bFsQbETskZISRzT+sUQAFQB8/KUFWGLcHYBoxlL
W+bAKiClVh5/YKnygcvIu82n25FlA8VyuQIOZd+oA99ileYcDpay3RzZhr8OtNH8juY+NqFQQzHX
VU0TLsjbT05Kp86QlY+n1nEYeakrTnuvrn+twTcurqdnq33yJDLdcUTCCcGvweSh1ENqSSu4KxFE
t1QvoEmyQkFZlT3Wwa5M+8ew0YHU3oMYy5ZJxFKRpxPNxjoyM8aMQlfsUrwdhVXJjwhHSqxpNgSS
hAip7GaRB32GDFBLrJsZEzXG4B7AuZUcAip6IA0QB2LhpJYIO/WTiKSXgqtzUx5dOe7b/u6W40q5
OGWt3k8oJf3LsIKWPIst/7AnwQV6uII5+8Hzu6icVfbh9Z7bge/4PwBoqG6ZTHfVtVZ0TBG2ySem
UE93yO6Fza4Q+iRrsBkcd02ixOXa/KJTdLO0TclyHMVJp8Lc5gTUtJwJz3d/iZgk0t/xCAFrM6Ir
MG03wFHdCp7n7qfYbN0W4wkaF6F7tTKh9asCh3raLd/YxwDGj6pjMOzeKcxZEWb/0ut7xZEU9Zwj
4BV5jT/nh1BSoY4xHr2xNXASi9VuaFL95S4UmjQKuIyh60DH/EcKH5OIdDDLgs54XK7jLwR1PwxC
zcsY/WMxNR02HlGpdv8B5WyLp3h/PGU9rGBV7E49SCutQZJRKy0lgogpLCcloluYaQI+P7yRs+Ae
/I8uXCepuosAonP/x8qD0UksFkNC6uskTnnMsBT3jJdywGbkVDhkDsRkq5diAVAP9iyL9gp4Ss24
2isx7YCrqUdlzS6HsdKyReVJvdjPrD3aNk+6TANXyioNJqhqIOZawti17s7ghjPopZmNaEJQ2jEx
zwZ8tDOgD23unYDADxBfXkMDavFmQtmGVD7/FZOJXaCI564+wERpkF728nJ7cWwpwWbJumOS8NlJ
KE7rss2m6V8EtMLBghowWsmN+kBsdYXmFmOV/i7EArXfLcNpNV7OVwVCz1XdnrC1HuhrYh7dDBxN
3Xk78ashTuUQI9oTAnZRk5Z4hmntlRMESiNBMtOXUCL1tbtp0ywGAHIJcvUztYoyUsvYPs0fSeer
BiOXMicPBjh4Qj4dcvGqA4c9lXw7P+ebM4wOE+Tel5CHgLbSKT1NptWzZenlE89Mq/nnxux+yEJV
xBZLLhxUiBaOxHQ38fkUIgmeLmRLUO2qxvZL8Xd4LO3vD4SjLaYHns3H0rSTrIW947XC5HMK4Vht
jnJxtPAqbGOG1RwxRVUY0n6ljq8XNj8MGXG7qZfPQ2VmNeRjh08yuSr34x2xD0Onjt+y2kO82HvE
TIofLJaTN3knKKektmKaD0fDt4L/SnVVRNPopSrvPWR3pL78JXT5o6kiRDABvMAKMiti6haST9/K
IDQSFhbUA2XgflP2S6t1rEy9WSZxfGw2pL++9xkkTOl946PTyUcIGFKX+xF7sca3wErq1SYXenyL
fvyfH96jsyeCnTncmcLdI7erlnIeEgKUUdMdpQY1Mp32Ry3F/1Bif2pIUp6Dtop4yYpyI1eKIkXw
WQ5IDnmfavs4xRm7ejc/i0KEsSZ1xBI0DkylaD5/UZ19Q+OqEz1pfa0gyTR7A9K49+dBz1oV4pp4
fAKwrfEmYrwUvqfVvjq67VCiY3NFp1Ov7M41/xsI3qTJgxWyoBpBIOXLefXa6EX8bZPqwtgY4DFJ
U6xKUfqIqIiVe7q0BTroNxN1gmiN0azjno1RvVrTv0oJTsp5Tqdsl/ShT4d8oW08CZA6rtx/Tndw
h90+T+yS0GO06yhqa8nO1n79dKst0Bmt72TeQzsvaLlKRKCPE5R/6Yo2HFUMJkq09zIQm6gzL5Bs
1sC9lmkiuF+PN5wGKPCalXkSocm7+JPUaSf0K/u4UuBUi6vlG72tORvEZFxA6nx6Yx2Uiaks4fI9
S0W/74c+G6NHJ4kLApjatVHA04fkDMnjnULwTsVjoWEK5zPr6BuvbR6ezC0OUTtsyOkMJRFi68NE
yvlZV7nbtW817GlSaFf0Esvi1ZbAnH6YzFuyKcxbUVqKTGyD7DsSta/EPh/9I6H0kGmA5BCzOdFv
Ca1LHBSI4oPPJCiut9O6Q0rKHUe36ax4pXjYRBXpMHSjjZ9Sj72nF4WnFLPz5kHfbZBT6FeqvTnB
g6b4wFdRoQEdxI4lVf5s+bgEQrd6psqoiT54Juj2lC4Uw3BKiSLvAcxB0kdFHpvba6P9tyi/39t5
0wf4iLHprKtkgZlv9qrzdzOo7sHUZ3b65f9xKZVBNnJOhrBunRiVQaOTfH8wpuCsh/jf2R01LRfZ
nTiDmvAXJGuaNCQYw4StZ6RdbdeADKHAGrtCRm8VZYuo+KlgQLtc6H2lDNTqqu3gx/JvmwY6pIaL
Y25hayAi53rR8KJX4q9lnx7CHjPb7Z3HWtQxbzxjue+ADj7Mbtz5NuGe5FuB5sgKZOYsBh6B5ORz
MZHnmwaW3+f8xN6v1teBGFf4ly5c6TOpouXWFc3novUi/9r6V+nQej259/jISgVkXdP9rT/G+OZS
pyPl7sQx0RzhdvO0/YbzIvGLB442ol7gYjA10MlALXuQtHQRwG2xappqkCiY3jullP4h0I2Dpwg3
oswz9RxAGHAflD6AwVNFvdbqE0NKIYd7MGAG2zkj0eIOXvMvvgF9g+H9o7KHLbl0wu+Lwo5RJPzW
ESJci8Pl9sPpaa1D9H6JovOsFQki9TL0hL9Zxw9BCjKGPwj1VOGg3hCy3Ligx2VRvSZmkfottA11
tkD8Drod0LLUkYZGaByJqagbp/Fr3T2wtkYVEDoThfVxSKJ3+FLR4X27gSfsJNHbkdXikNMgoV7b
1F2NT+xDG4BcLTucpMUCMjRpEDHeUC9b3+/dn8leyvLmG0obyb51E6NCoz4eeTjGTd2UBDK3sMeJ
g6euEvYmH16cs0SlRHv5iFaPI7ZTGrmv950nllDhxjDQc2yeARhirZSZDVRPWdP1FfmE6llKEH/l
UheNpZJzfYhtTZqi+3SpLpjHAayGqbT6Sk/JZZitSrZSft3bKTFb+9OEy1vHLBmFwlMX8clqlNp8
cpret60YouKiH8mGw1nJPxhWR7SysxlSqNCaUkPJ66svo/b9BEa+5p/en+8Yfj+RuRqOqZZ1abcF
sqfqppw5BSOskRtWPF9W2hkMCTZCHg9R30T2zxF5/rb3iw/FYQNpcoYu33PRmckrFFdwSK5RtTfP
c80ou6Vb274z5rUkIE3FszN1TiduM/pJWuOSl+Zuedo3Rjj68B0kyQdCnfM94EVSl/TIz65EDAjB
hx9SYgkTjmzbGlTmuWfRl0zVKd77MLDwYeoXa9eDIzCRY6X/TxIP8Tz9C9h6ZrUTa2hZYqPvGfGd
Tgb1bV7ttdojPYb57tOC1fW2rJKCmEL3T0umINZ0Ajbsc+sCs9KPbNihWHM1HuLasFSOeszSun0+
XWe629Oc+ku/HeG0C5CBTjfj+46xJ048KHJ77MAFtDgp7BmNxBO4BksC9e30RAZ8xnMcCzXR1Jui
+PyRk+JvcdgiQ6EbLl0sUP0/W2nRMekePzCQSyCVf1GBxxmsiC3VYXnmYZkTtelJ30vW3Zm3oxVV
VIXP7WXQ9/1m5+4Hc5BlDVrL0I3oo/KkGC7W8f0xfDEQfDPF5kOWFDSDZgQxG4lL2xSR9G3mlFq8
AsZf7oEmY5xHTbCQ5uSacMCadO41ADJaK9Q3ZUVPYKgy9hH7ciVZYUoVrzsBAmLKB929hJdcNHiF
rox601cEyQp9I2ShdETxSX8gM80CG2k2I8+BMrpRCy5lN2laI3uPA2vT3WsrH+6ob2Z6vdOYXEPG
7sqO6X7SC1Ptr8vLKYMjoFUWF5if2rq8ZQynajr2MPRvKPDVt09+v93rTldxRTRBGU8933PVIxgk
wua5+bYlSLmmZKG1u7OXi9VoGCXBkmIo6/2w0XPraUMNUKrHDvtayPFHQPYCkmKWXbcw3S1jEc48
MGPC5s9WtTuqrWSyKsZzawNf83V2gYHAxWGQB4o8rVygIZF5Zlu5YzLgNujAbfeZNt5PmaqJ+CAd
rKUsQF4aNhswFFDLWU2TrOqjsO4zffQBVmXYWoib5Dl+yeYiYpUMVTh8qpx9WMjtV3iEr+12Tqm2
B/bmitgGEMsqjf392Ya6gU1kQDumTnmt38GgmKXUHhFVk161sbFeL8YPCBPRvp9uICSeoGyhmL/c
KGasDsKqJ6pj2Uz2EhJzeM6gx2cTmTjq05YmnX9cXE63wVQFOx+nhQlHyLhbWx8rnbp7+p+I1/YV
bk34YKOptvVYNpf8JpEsbY+SI69AdQii2imYV64eLRiFtcOBvvTk6ZsrDqWNMOejbR+Ot3kcxcPB
QsHtixM3RAe2xS+dux1p+90DX3lE5RpBqkWKm18XsN7GRQc6ewr/tTYaJxYwvx5mcEM1A+AWlMLX
U1whHziqgC5487tK9FkZstOP93OyFuhUtI1AMUq2W4gRfwujhgl3sGrFANTUN4cuTlazvmpQy24q
+phaZopznJ91/FAmlrEP+hJ+KzOkxfNKj6S82wZWCMNmug5GZQin/8hkgznQXfHNz/tIwp3AeOmr
kounUsowzFwYw4+ZL+W16MGjKGt4eBzOaDm0XgrA+IfUmUbzeoqn00Z9sT4hmqYtfYQ9SZGKWzus
AYB7ypRHBN4WRnaZJ97xw2F6zfe/cfbFPiP0M+GCzjG7h0viQEtbqtXUHFl8EjE1JYHF4T67+pJc
LZLbIDPj4IQDvVCSvmhTEOSRZQXD15MTU315JkL6pe+gagKTiG9ISdMnPV5fHx+zCsHm2IyKWfxF
nSMgwT/qfT9RX4mZH7IWNEBfSx5Pp5cX+G1jy7lCugGOFzxBUanq9oQLYh/q5INpbq5jADNKlFdR
D8zcRQPaPY2zvII7j9hqP5nO96zftOo6ojHtUelnA7JZ61DZZrwew13rle6+x8fI36b/uDc31ZA3
MLsgc5iYbC4030f3NOvfpyRi9W4RIcDkzUb0uTuy3t9oX02meiO0s0h/Ds9gXHx1ShJ+RNocBVvB
xEDPt8t5Z3cv5gegwuxwuSJll+7Knv6ECNATJv3fS26TRISgPXxo/QzUYSyEd/SQt2yZEjSRUKgk
7kKXZKmb1kKzkVKsPVl/9gkl/58IqGzRgwkh1sPN33mKOe+icNkdrd98FclH39Z9GhW9oWOYljn9
uPZXHnSpufVGxqhQ0MJwL6Qi1pW8lLSwGMjy0UWqNX3rG5mErepEG4zS/wZP5r9BknmErVjgyw9n
LwXn2QTbP7EqBWgL2fxRJt9O6LMsAxdzVE8OVmztJbN0w89lKNv6YCNfAPmK0SSuK0ILPrdduhZw
AY5QUT31yl6iMDVB52Ig+VJ25AKk9WtGi0VU0Yc/7RT5h4U+QcnvUPIYzxG3KSr6kdFRnp/sr1g3
VAC9kLTnMCEEkaVQnCOwi7cR83tziu0sQzz7k4BmDJ76xOQBRS6vkZCwXsr9C+5qwJfynNGSKgib
8XfGwURLDNsBUrCPmPx/G6sSxIVaRITEu9uV+2QSKPgL+UkCWD5FfZPzWZ6Tg1fcUlJ4mKdnttjT
7P6YltMo9YFXnaK0gy/hfyZyECb4R1pykNGgzueAvGLQCGudhTZVW9JQwVrZq7FMeAwWbBqORqkH
2pZyWfaIxZcRYbchBrIjsSA1W0RWV0rkmXpVbe1pDfGAdhXwLSq33KEsG4fW/F1aycEv/+bFEgPU
TGJ1X15Dq1M0NaLmTmA389samEpZzOmejkNftldsRUf1eis9XyAFAANV4YV9BoK3JKOjV5azEl2P
OdLV4/GVO9mAPZQReXSXbBAqe9r3cGhAThQA8me+J8V0njJqTYTAJXKE+KyfaEpgQ5M3Dl2NMWwV
DWWa4YQiKRKC32yNe91E2upqeqEmT8QGbw==
`protect end_protected
