��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��33�z_�`�f����EW^7"q5���K��Ҋ���CU���w����=G&�ʉ״Tĕh�{%�E��ڀn[ɥ�'S0abx/����z�K40"��bYʑv����(��C�)�'.��8AIH#Q�|��H�Ǭ�Y �s@�_u�-����A�]��
DL��T��6b7���h��,�x*uv)=�R[��p�>�gr�N�a�sE��P#Wʍ�vfsr��!�߇?#:3N@I��D������Zz����%V�GE���.�$�����t	,V6�ʹA��Mn�(��<'�3:u$�S�A��;�{�9^�L��+�PV�f�����N�?K��|�}�����h�U�(?_!��dvc��-!ԇ�
t\�@���K�is&]@C� *����f���tNZ��i1o����m�ZQKڋ���4�Hoq��/� ;�3��/�'�jju����=���c�ۧ��:d�@���]j��Q!Zk���~Ǚ a�=]�^�ڻ��$)��ans%��ƫ
_�Y���ft�;����c�L1*�h{n�ڰv����=����Z'�bDI�i"F�q����U���/L�xY-ĺ��g���7� �Q(�3p�$g^��/�|Oӛ�;ߐ�Y�%=��M
:�T>e�:?��y�I�h+�7��x7� O�EFc(�gT���������8t$BZZ%���K�+wg��R�w����HȬ�{f�(���Pe1ۓxao��nj�ͯo�j�+���@~�����8�[Е�2@B�����05ڕ�}��hQ+����&~��%th4��/ �a�tS��~�I3��1[��i�|��d��3�{Ö?h�Aޔ%������ͷ�\�ܤ����1\� S;^z�L�ĳ�f9^M�,�h��L�)��<�&��4���W�ز�v�7 �"@t�O��d�#�uy.�]h�'�Yp�l���W�ҷV��()C��t���լj��t��,次�ee�;�$�s� /�����\�U�bU3z�z/\���
�[;M�H��i�a"���m�0/p �["^�lO]Ef�t@̧��Qr����a/KXn/�ܬ�vm��D����4��fs�^	��>ۖ43���l�GĿy#��h1��8!��Ŏ�����$o�ջa�@7��3$+@��z��ܺ_B�su�� v���s�t]&����7�v2�͇Ŕ�ez�S���,�y�V�b��,Z�G���+R���xO����5(�G\|��g���4�5��˒@�U(S��45���Y�����^.��I��CZ���V%p(w^�G� Y�}�z��q�΂aa��X)�H2�de�ŋ��ӵ�����֣�-IPGq?f$��W�GnR@�?hR�?�H�yj�3`$��.C�^ƣ������"Hy�!�tگ�S���j����^��@��x��u��cm�H������vE�5)P��*轵�/64�p���l���OIx�e��5k
�$�I���z5h�v�L���EkzF��g��'�Vs���r�Up��A
\tzpW,����ǚ��!彽~,:��ӑP���?��}x�YOxW��a�;��Q(�e�c��P���X��x�n-��vCѧ4��^��G���7f��� ��V�:��Ly"D���/aX���5'n�NL�笩E>U:��رWA�֥w�.��\=�3�d���eAgrX���a���#Z%K��1j�{$s"]�Z|�� T�x��i��'�J���Ջ����������A\�G�q�����B����T����գ�=bδ��)w6S�t���lm]ԣ��,[�lAǁ3�l��8^'9ȡ�qS�/Fj$��,��o�,��ڬ��m�6�%!w�9�r�%f����}6�e2#�v�iJ%K���	8��� �R*��^X �迎뢑��1J(7������%o}����hH��������pwA�\{L���0
z~����B��]�|��'@�=#{fڦD�S�!����o��eu��[6���j��aڤ���K�c�ئ*5,�lV �@��r����2s?��J��t��>���L�|�9��$�9L�*�=YF���!]ζ��̄��|Jk�m���ˤ�2�P6[Ń�2�>!"w;�J���n�,�4���$ 2z��֟W�=0
Ą��o�'z&Ь���a��k�i �n1\*�Tdv5��Gݝ���'$61���Cna*���vR���QyU[�L�k:[O��	[ ����(�$&�e�2+J�9��N�x�0s
=����׽o���0�<�Ex�yYAj?�I{{W��&�j{�0��o1*}|<!lJK=A�aq-�*�� 9{�&�P��j����i�����XO��+���_0�	k���<)+����%t=�t�����_Ȼ�;_����aE=��6i��L��kf�[�{_�z�.�h3W�d����"A�jK��z�x����H?\	ڎ�V�E|��'(��	ְp��&Ӡ#�,�q؝G2������U��hUQ�Y�a�[Y�F������G�<}����#/�>nS6gn�ڠ_��E
��(���ӂl?�s�1����]D�3���d+��Om�9?��gIƋ	\Ŝ'�ٿcI���(ns|R� �ci^�%]�)n�%�&]^�If�'��U�b5�q�bnq�˟-���H�E�;3��!⽔�<5������'�ȶ����q�Wӻ(>�}d�� Z�U;���5�q���Oٯ�$�YP����𙟏[$
͗�<U�Cx�y�k�J�+r��ꐞ��)fn(�l�l�a�tR{h^��������czr{Y��"{<c�&8&~�)�f񤚠e,�35��>�ۄ�|�g�Y�Y~�x��ƞ��x)/+�/����9������~�՛t#�����W�nOk�no��B��)�S��RUp/�'T`@���������靾NJҽ/\m	?�p��
�/��D寲Ht@�'�]x���;VY��娋9�'���W�1��?�Y�-��� U�0�����k!A �X�xD�"�(��(w,����XR������̢JA�P�O�uI�E��1������Hz����Qm5af8W� (�y��
��Q"���5��Hok�����6�e�R5�U實��7��W�gG�A\��O,(��X�����2*~1--"в;����D������z�<Oz�;��v�Bˢ-���z�/.����M5��D�`�A~R��ˡ���&�C3������wH�:��+�+��qoX�[ܪ�	�J�_ܰ��
�.D���Re6���!��7�U/3;��hT�qp�"������-e�c���Ò���F�_�<������O����-�刽4=K������cAw`e�N/��Hq|W����(�@Mg	�� ,a7�tugP���A.�x݇I}�^�y!�u:z� ߻�h��,���UeO��<Xj�î�����[nX5�