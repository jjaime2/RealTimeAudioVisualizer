��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊�{�_1#N��	�Iy�(V�+f��q�>�,���ٵ���k�2�'y�%������7G:;���0�ygվ�&}{4�6Z�hi��T���-B���.h��� �Y㷄t`���@l���"2��i�_<}#�c�Ęٳ����6f���pe~r?`U>��*�lphwB�G��av�WG�I�ܩU�ʊ��2S��/4fyT�vF�i�_ /�c�WG�a�*�\�!}
T��<]�#Wp_8���ũ`-�ݟȑ��规��[�ձ�g�sE������Lq�E�LdO;����.^(Q���ٿ	�X�V�5M=��E�w���/�jF��w��cZg�Kx��iv[gA��X�#��C��/� z���.[��F��PxL�o���}�W��v�I����S(�}�>`���,x��;����5���"ֹӱ3���[
���O2^�E��&8�|-�`{���Z����8��O\W����n�RQa�]H��Q=[���,�	���~�����ZEؗ�%	D)e�~���C��C���h�p�t�"M=㫧���n�e�Qub����}��F�P>;��MZh�U?L�-�|�V�p��x��?ҿ0@�A�炿N��f���aG�>�D���A�X���٤�ܹ������K|���(Ad��dO�����U�'�G�ހ2I���ݗSjN �%d=�����3e��i�_�����K�>���?�?����r�Ĥ-a�/h��^�%���ш��|i��D"�I\W�]YBe�g2�I�R.���G'�:����������5.]Ĵ�"���^��Zކ��9KDx�����y��P�`��mթ�H�V�-Sv�4�$���"2�r�~���wkDi	��G#ۺ"%�k����!KP�3�E��y;ţL��D��<�l�9��PR��ͣ��!��DO̳4L�Z&Vӓ�C������DI�w��1z��yN���ӛycu���D[�2��؄�����K�GT/&ب���Z�D@8"��|�=m�E&~�=�cs�6��Rm�߂��+n&�܎><|	R�t$g�N�p]-�H�3g��З��s���+���X9(&��_��}�V<�Q��=-m��
�p�RͰ�Y�$�mƳĄ��SG⼦���rD�f9���֯9F���BE� �l�ٔ�p_��2�tgw���b��4��3�� T��Z����6��#�b1�����&�r��f�,G��'��J�
�Q�4�(��M"	�|b�H�e���J���ߩ��������ߡ������;{w ��#y*9fO���O�L7�>?�/r��&��9
!±��YD���ċJ2�F3(I��t��:���]TgR�2,�{=�h�W��W�Z��˱.���K*������*?Μ�l���گV7M�Q�@D�y�C�=Bc'98�J��#q���Z2�d�st���Ds�P�ؓP�y�$�
п|}�<ј#z��V������3��=��z �U��
xbO1c�L��s�QΓ[q����
�-��ud݉7ujAS�(oq��U�	�/+���ł���(u����It�Y���{7	G�p�˨!e��c���Mf0�T0��C��P�|�/�d�X��^Ih��OH;h�-�� n���>uůXܢ��V�M= �W���f����gp �^&YK�}��gQ��gX�n �E᧋��:wd!��?|9�!pQ����oz�'s����a�|��ho��; 	�CDp���c�1�\��v�D�L$0EK����S}3�a ����,�!Q>��<�t������ˠ\�g1$��C�\&U�"�w�hM��="3`U؈c��UM�6�A@#_��,�&�6	�.�UG�Q���;���e�NJt��1��c�B<�1m�N�^r<�0\�˩��g�?A�N6�������?dB�K��>4t�R�ũ��"���V׽���V�O����e�¢z�K��qV�H��z�	�����áx�6i�֎@�m�|�w��*�UP[���_`��J���ڐ�R<�,�s�K��O������j|-۸-cg倫^�A���9qէ?]A�@~��&<��oV��̦|85�5=#8���� �R�s����\��G�t���o(������T�v��7��F��a���?b,6�U꿑��Ù��X)(%z����&0�J3�-6���ߢo�	n�#�r�<����B� Gu�ToWb`F�)jJu<'�bkx���k�N�/lj ��I��Y�
7xI��Ġ�Ü�	��Jy����|��=�C|��zM��?VvqB�p%�G�����S�aVp
�]-��D�;	y���	��1����~|$u�����#��\����h�gsM'È�*�[B����)�Cx+��������gX��d���}��w]j�H�õ9�A�U�f�\�SވiˮO>-��.��j����7ӽt,s�������3��i6��֔��^JW� ��J���>��3�6u��S�~ѣ��K-)��@�[cI3��f�u�0,��K3�M�tݘ��B��԰�����t�uP�����I���a����#���o4�1�6������+�7�3`{����.L*��	���fL�Ǜ6�E�#�b����B��c�|�F0}�d$ s��ZT�;܏
z~�)o�Ky��̸����Z�FY��c�[�'�
@��w�|�������;�s�����о�Bө�+L��0���^�Y��9�V��G9��򽖈��(IT9}N㸙=�����60R_�
1*�I =�.��<�BU���gW'4E���
��=PviR
R�Oy��Ls�B�xo+�]`#�YrS�ry��q�9Z�X�G�K>��(�E�:��B����:�Fn�Ȋ�$ѹ:��я��Z�a��u�����%�u����}�GW ���s��R~�