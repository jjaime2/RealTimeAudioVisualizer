��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ���l�$�'�Z���u��E�a ��B'v/�γݩ%5=F�7z�N?ysV�k�b#!sI[-~�G�m��]v��G��&��qx���m/�H�w��V����f�Զ�vp��B��\6�Ads�-����jfc`�kQ:�k�ɭ�|��&Υ�B��n�R3l=���]�_���Ro���*s0��|Ft�m
D�e4,�t�N.��a�˽�T'�C<`�e����E(�!$r�)��}�����3j3Rċ����7@�(��zmt)�`��L���Ì���j�LWS�g�K=.����)	�,x@D:���y�!_�/-3m�o1�ʱt�ŏ�z�'���A��@k�#Nl�pͼp���I�f
�KcF\�2_�SY���'_�B�\�ݩd�t�:��q �c�m�i�B,��K��ɖ��	2��ƃŏ�71����)���Y�(3=P�=P���Ɨ8�l�^�ݓ�?,��Ұ�=��H�/3��-'X�=�Xו���L�K�nlo�N]���zY�"U~z��b�B�?�yD��I�ӜU�hg�W����W�}��1w��q�i2`�o��_H"��Cq`���i<���l��"��
��룱�k{n�	��E�s��O*d�H�s��/_�{`E�E�nQ����Eq1��&�4\�橕�`�/���tl��]^6(G`��KT#{=�L��5�BN.�7㭴�̨j��ߢ&[^�U,hOV'%�4b�Y�1�~9�Iqs6J��P=��=���x��~����i��	+1Պ�2��*OhC+M!:���z�0��j{���x1��Ց���o���EJm��CJ�~�����$T�(�A�����R��.�I����;�]_�e�u@��DT �-�j�=�|�����M{����65���bW�,�K���s� �tǼ��o�AE��"XX(H���Quq�3��0��n�[1C���%�!���(�8�N�ӻO�����BX�w	[Ǐ�.�)�?3�H�mz>yo���6h�6D���JmV�?9�q$KBP�Z����X��d�sC7�ι0��V����l��|	}%l���]nS���_6.E��k��+T{6�:�v�:~C�ء��ak]:���������˃���B��,)5̕9�)��ꑤ�W��w���5l��n��+���(=wL��bd��@m�+���COs_b`_)�D��2lK�Or�:,x�C����O���w�W���)à!�$��M�U��-�l�� ��tn���+��rtl�d�|�m�G7�.-(uL@Fo�>ـ7��5&N�;�*i��b��7�Lv=���&����[�����4�z�',�oA��xA���={R��sY>�G5�2��w�s��x,�n�r�$������Jh�ɥE���˄g��3Dh�L3wȷ��)6���� ������,&�����d2����6�.�. ?/=U�=���֮H#�f]�����XiXUBL�-!ǣ���h��ó.�W���}<%^�<��(K�����g/����(!$�%�a�*?�F��.e��gL�dF��uN����}AB�
�S$�d#���h�7db-���7�o�Sb�^+��������Φ�\�zA�o�H)7��u �tc��+�������k���������lD{��x�{�)@x*\�kK՜-ɞӦ3_"��؅�P��F�M�Z7}����G�|�J�j�U�xn�l�Zc��MO^l�.t�GU{��_�4B��]v��ς��yu1�{�^[TOMd�Ϗ�ey�˱��0$�?����k���}_����wV��Ɣp��Cʌ\��n�9�OѴ�dp�7�L(�j��ZQй�04�i_�mWu�'	��vT�/%�2���M��݉S'�����De��	��=�2�� .�����z�1&6$a�X����(�ZN�y�=���er9����-y��-}�����3!�)����;�d�LA/�<��1̻r�����1$܄�WSf�Q�(ޭ�{�U���0表@~/��#3E�a� �3�\�֠e6��2'L��� �H�yvo0��	�]�$�2q�ıfQ���=Yl�������c�˕^��r?U��d9�p��� �+h�>=���vi�m��*��,w=ˉ� ���I�}����副lZ�f�qTq�h$��aKd&�!�<�JVV���ݷ���
?��2R�T��k^�Dԣ�C�9��뒚�#)������b�
���O�����k�'�����>i�\\��ҡ�M�J�f�1^������J�B>7w-�uX�UG��W�9��N7�`*�A�%h��Tj=Tw��ZQ D��.�|�EO��a�6F��;��|����W1��-k�Ť������K33��w�8��6�ٓͅ�vEq���&3�+#$�_%��lu��-[�/cB0a>-�c����Jq�U�#�2�	�O"�>��>�z$�6��tݮC�����bz�d�KTm�L`%
MA5*��BХ�l��Y`�F�p�Of
!�we����}��wM7S5b[2�G�?#��kwt�d{*��%��(��͉<�V���vN��<Ԫ���$^�|��Yv�0,�3����{e����g�Xo6�+�r��\ė[���4�)�� M"�'>lA��v��:�����n��W�K��n6gQ�MJ[7̗�z=����1�#�����`�g�n�hҾN]�m:�J�#Pm4!��Gw��`gu��0M�� ��t,�K�2�r'ޙ��b�;/�����=���YI�5I>�ۙvU���6�-�j�>O��q��~�Rb�q�T"���Aē����$�f���������*�%!(��sV�4&@�7����`Z/����5�l�d����5�͏
G1JB׼x����P��h�nćϴ0{;Q�ޢ��}���]�F������_�]����c�S���>��Δ)d1����p&#�b5K{!�to��;�1�տ��v�� P w�v��VS�x�LE��UX ���rL���,�� <��^�B���)��?��%�Z�]��0�	���嶄S��4-k!*��FvM`������.���ެ��������4S!ђ��L荊x��(ӆ�IV߸��]����f!�(E�q�Fv#]�f^(3��L�9��ը�vu��7���m��o�������� 7�Ӽt��Vړ�A/;��ޣ����?�� #��@tʿ�d�i(h�V���?�$�&��ݾ��w(�[r	t%v����S��1h�.���rGԻ�,E�oJ0�Z]�J�/TX "I*������k�Щ4su{c@t���G�j>������b��;�Z���j���'�`E���(���w_U@߭4�x�^���za�&�5g~�_�i&�O5�e�ӿ��V<U�E������P�|�[V�>��Mw���*z�&?\-�����E�9d!��ب�MS�:Γse�ͺX|��z�ELa	 ����4��H�ת�A�"9�|�D�D��B�FqV`�*��5j���E��DGJ`��YV4 -ߥ"?��3c�����\^	�&�zw҈5Kt �`z=�1Q��0r%�y�ް���wJ�3�W�J5��bm��k"�Qlc o�Yby(2b�"�!�vM��ݾ�f�v�w�7��Ѕ���gD?��c�^P�}x�]��Ep���.��4�%p ��'L��ڭ�'T�g	q.�%23�+�1d;(_x"��`:���l�})��~[F�4�_1n%þ�H��#�u/ᮣ\2<G:�&��^�r�@X{���  \�;\y�^o��<������4̀k`�)����drM�V��8z"�.4���ÌRڇLL��G�qD��A�c��8δ;�+�<j��o肛����u���$��B<��6���j�<|L�����%Ct�[Nj�@�9ų�m+?�N�▍ '�� 6��I�!7�}|��e$*@!�2��h(�a��jM63��ﬠKY!Q-�X��`���3��^0U�~�N���9E9Z,�K>�	��{����ɳ�r�A�VTtx;H�R��cf3������y`c��h�ə�K�C�C��e�$��Ð0<�Rb �9µ�8JC�gv��,񨻊��PRm��1�?U��Qu���"S�d��sE���z��;��醇+(�R�����5C�ߜ�~���������N �5*��Xc���Re�0�����7��|*s����lT�@���6�Q�<h0�0��<�Ζদ���/����T�����5q��4������|>:�����$����/g�+�6Y�T�̰?$����(����1]Y��΃�����M��]�����j���'m�^"�7TrrW��B�QE�\�֫� ��Tb!L����'��3�)�#�7Е�Ϩ�ޤ	w3�hc&>��R���T���}��t]���4v�0�mV�ґ7�_�R�,����=>d�R��à8a�:���`R �]�`Ky��o�_��4$�L�-�`r.)�ݖ~�^�/��N��P.nO8"�q-��I� 0�&��ɠuj ��N� 7s�Ϡ(E�a��q&�^D~���>�����Vn�τ�'ɲ�-�R�+NSC�K4'�\�$g�H�;�2Ӣљ�WUN�dq��)�H5B1��抜� UajY NB���JiT�(�jG�����(o�j�k]5�*�jGQ@"��h�嵱Y�1���L���B�4��R�)�tm�E���tT\�ꅺ����BX�����$��Nl���� �~?���A9�W|���;� ҅|�t�����w۞:E�x؄0i%H8l��B�����6��N_>��h����le-�j Uu�O��Z���c��	u���4$������Zb�����.~������[ҧ�}�[����������wQ����-��Ot�R&Y
@q9���~�>�<����'��ί{Ȋ����%�r��"IBA����m�ϳB�ƞhx`ؓLz�R6[I�T��)��KM��3�&�g��6�W6Ә-���.�13�V9���0!��ڭ�|�Y���*&ٔ���$���fP�UՍ^����ά,�6�[,�*�d� j=v��-��]�U"��h S����㊍�"�x��3NҤ�RM��������WՔ�һ:����	E������O�6�,h�;�Q�09�^P]WI8�-yV��q��*�-��Pu��Yq)�Y8�l�;(�r�R���u�j�/��Ռɒ_�+�O7^[8&f>�~�i5�̀�	�?A���j�G�qY3dA��`_s°ZONA�؞�ݶI!6�lS3��%��RC��:[�s�_�}8fs��lq��엺�d��J[?D�b��3՝.k��%��ĥ>���yf&�n�e�IfD�|���z�³c1I�h�{.@\�%�+,���h����7:&�,N��:���fV��Q��
f,��kJ�'�~�75z�~%�7Pju�ȕ�qqR�̽@i��Ơ ,hf�s���M�yt��I)��.����_�z�����[���k/�t��-����E�c�,<����h �&ָ�(@���;�T]`VRx͂IR욬_��a{���H�o�U���ds1C`;�nm'���V����w��K��� Z������"��jxW$�LOg��I�>��=c��W�l�j��=�����6�4i����t=�Gׄ��|E��B8B׮�!j�S�o6�Dp&��[h����3��t�"oZ\�jV����y�jQ'4���M���������p��W9e����A�'y� ����դO�0���x�ɩŧe<0�FZ��s�)��OU%���I�FX
4��H�W��s��`������]5i�D��Qw�&6�G�4-�	�|hP����{׬�gd��^/��U	r���؉�f�h�S��'@�Ea�����(��H�L�kD�/v#ٺ���[ʗ�%	�8�����lֲ ��P;a��&��y�z�S�M�bj��q��
u �0�i�Ȅ��'x�l�]E���̮=q�C�Ԩ���k��0w�	6�m��u�J�v�R���s���i�O[�
yf�!ˠ	��?�b�[/�i`~�t^'hL����ے��Y�f�������g���T��/MQlp2�<v�.f}�Ie��@i��ڄ��]ಸ5@vȔmb����.r���h����D\1N{��p&�{�|>.�:���n��%ܼwֽ�l^�Q�s�s�c�'+6]k�m����ZB���<�F\�$cC�#?�
�ym�a#׮dG�.l%�	Kt��a�����?�X��	��_�?��B�C����i-�ɚsiR�+����O.W;\�}����v�1$ º�I�ؒ���]h�7��rf�y�PL�� �
<焫|�TI��g���� ����f����=g�������^�1'U�Yƕ�*�P8xm�M��� ��x�����S�&��)�}la�nY#�b2�BtJbIu�(�����K@�f,m�Mq99�WX<��Z�{	�{6i\�D��.l�d��!�=��ġ1��R7�?rٗ�o��d�
/o������3��b*5ԆZ�q�8���ؗa��诵Y�&�U���R�\���VEK�G��i�I�fe�*l�m���d�i0�fH�T�0�N!Hi{rN�&�FÕ]S�B�_�i� u5�n��SToiq�ؚ�M��F˪�+=N7f�0-I��0T�=%6���ԧ�ۓ�Ɏ�p����@����I�U�g�A�,�#�y��PϾ�AƄ�~_n�~W���4���YoW�Jt�@�Ħ��P��>�}������؇-�Y?chE��JB��*��>m��*'j��YXю���s�lޓ���'#�En�BI��l���vYX!�W�"{�{�R7��s����w?z[���J8E�5��IJ��t������ʠ�n����#ʞ(�v�0�E�����b��\F#a=����x��[)�h�fSP���V���c6�ng_m�1�<��`���-���h��kN�󭤗��{��`A�w�v{���)��Ñ_2�]j���゗�7���ٔ��� ��&2W�l�OCqZs1X2|�f��X�
�����p`O|�	���C����a����7�g ��V ڛ�����e�'Q0z&��b	v�Ѝܲu(�1g��iK�$��V0T_8��v�M�D�X��Ĩ���,S�m�>�`�onsE��Pl�7֟�}���n)�'�-�-s_�qB��тƻu6��h���|�鹄��/i��=�hx���&��yO5S�:����{nX��;;!�x�#��j��A_�����6���O� ��Y���j�9.PuźC��ǻ�W����ռg���s7/��Fn`����EY���5|��F/r�������Ƕ�5YS��P��s�R����h[G������=��Y�� ��I����k�>�;����D�1U��"��~^���G�/��l����T���ʹQNY�����I+ Y'Z�5��q��f�{��眖��xZiX-�0�O/�P�ʞ�B�[���r^I!��S��҅�� >9e�����O�\U��hN2(�E<�g����6兔��Z:��A8rjkx;�P滰H݇d��6�6Zڈ�?��c&��[^���H�.lM�
�����}Xs�2�c���������~t�V�(� ��B��`�Q�:!M���"���8U��@i	��h��/;�Y�W�S�?�GrV;�)���|��4tZI3H��.����pK׮ր ��ˆ E1y�qޯ5�1,���yb��V�v�E���%x���`^x�9�z�b�3Jj�j��K�q���w��G�Kf� r��o%�BK�6Rf�e"�~��v���wMj�ubC�Bfb�н���j!�s���h!�C�`g�OΥ}���e��YK����s�+b�d�Fh!��k�u�0��~D�_̻C�2z�0�Ƀ��Ϟ�	`~H�PɜYz��D��_�\6�.Y>9;\�=�X��vG�T�摤[X*-c-��3�`E&� �[x���*�gE�Up�V�)K�Mps1��un��TY�:n�>
Z�Q���K{�4��]\����� j��O�WQG	M��G2��@��0>p`�)`+�0�I���^4،�^��-�XOn0k�A��e�+��p��h�苁�;���������J��������W�G�u���Q�����*�Ѽ������IZE��8��̒���.�)�J
��n���g�{j��Ͱ��<�r�M[xfN"���X����4���.1��_Fu�������ǥ��d=�a�T�=O���K�C���Q��ޘ�����'�d��o���÷_-�@	a?�ۍ�Q�D2�*�\Ea�����N0 �@�=���ۿ$mr�yJ0S15bxPv*&�](1�j�f��Ƿ�.�>�ƛo�tS�z[{,�$�3���FT�M���� v��e/�cJ����翹C������b�E]�VM*�M�2;Us^���&����}���
��m(Mh �v���v�2��`0%��5�F�I��Jb�W���G�vQ�c�)�C��D�~H�K3���d�k�i1���9u��nw�"�٥v�d?�����N>*WM~�x���o_�E�������ɻ잶�5�ǐ��l�)���r{{~�e�s�(e�ġ5�KB�p�֍��YEf	�[�?FD��A����r�K��]��3X�}x�M�q&��Q��kC6,�`�-�k�g���>�IE�/��g�Sٞg�Ĵ��5���줚m�hk%��w�LJ14�)E�h�RA�iq��ax4P�`��"��Z�rA��Y��Ч���i�с]�d~�y��U�H6��FB��NH((1D�}��F�nfc"u�0�Ὕ�B��k�9�d��ʄ(H7��w.^�/]��R�C�0y�y��&J��~�v��iv��-��c�{�ͻc.8�s|�5~Rm�t�$��}�e���ڎ�a'\�wUxp�i$�y����^#�Ȋch�q��'�?G\�y��]�]6g����tf�K^��+�8W̝y�/�L���f��(}�������l�h��m]d��h����A���uT���\�=�m�"Zc(4�^饸<���:�P�Sv��W���i�l�����sC����4�Ĝs�L�[�-�Ԥ�n-�q[��?��׎4�[@��%�Զ<�H�:MW�X<�|J�����%���~�GMnܧ±G�+X�R�$���h��o�8&��,)�J��B������ |��ŷo�Ҕ�`��L<�6b�R�'O�,km|�Wn�ao�����&���ߕ���]��*/�2�Pi��R
����{����]!7�Ll7n��Ye
��]��Z]}��c��ހ���/K�G=�Ə�<.�����f.�&-aD�����,�S:,���������׿����h�}���ޙԏ�ղOj8vGQ�\�po�@\�Hs�<�xY�C����ܓ��8o,���FsD���W��ʷ<G,S��L�I	b<J�	
x!�W6�Xo~R��k}��e�[���0�<�6��+�����]�=+v�i4�!h�S�it�G2��8��a���2?�;����3a�U�Z��T�~w����{B,�,f_U���VO�#������[s7JĒ�R�_�����_f�٩�<Q?[����R����=Ё�L��%���)N�L�`=�SNW��Jx"�*�3At�����̟iҨ�b6�@��!HXI>9���Q���	Hz���Y0ꌨf
C�t��Gs��x�d��b����79��-gDR��JL�$L�f�hcD*�E�Jq�E�2s�-����M����_)a�x)T;�b�ĩ]hf/����ϊe(��`�vT���>�j*&c����\�j9ۤq{�����6��H�&����pI�3yz�B�J���o	�rT�����v�r� M��F苀��K 95�;�z�t=��j��
���Ń��ˍ�����1AL`�S�.?�#W�+�����9�����ah+� ֲ)���s����~⏎S/�� aWV���ـ�ɺڗ��&	���3r-��QϿ(�J���LS>�@*R�z��0���`0�sk�s��a1�
�[����w��M)�� ��0�ׄ��HI���Uz�	��ļQ�A+d�/�alCeղ���>���z��O?�Ի��Ha��E�("��GN���<~�f��RL��Ӛ��(���#����d�z����B����(��,�����ܷJ���<�j�����x�+9��6Ӷ�W̙w��k�m����'�VުR����G,�C_r$ѧ�s���uO�jx��$��c�?)S�#�ʞz�i�^\����0�ZγQ.?�6N=i7�Os��sp���+��]�аq�u����⪺OV	�b6}��[a#�>j]�H#��b��@u�A)�f��	��=n���E�r<P�x}������2��'���ɗ���% �|Bɯ|}���:�! n ���=8W[FK���V�n��~�n��MM�
�P�w�w�qU@��B�
j����
Y����!Xր���^�2PXq��=(	�[���aY(x<����P�'
����#9��ЇY/\�⑚P�����l��k�8)����< }H\4��O�I،K����Riv����!����1EMU���W��O��_9� ���Yx_�,^	������j:�_F-��1�B<&����,�9�B5$���4d�R�$� p^aj/7��+�w�g���4N���Fഄ(��Pi(�Rh��
�����PY?�Dk��&���1�Z&����O(]w��m����"�Y�X�\�h��3�aD��|��LU�'��[����vPF�Cku����e���w����+��Q8-�96�n�CV`�5��:��)���e��4ؗ���7]\Z�w��2��(�B3� C}� '����A��-֪�Nk�a�;�s���,�u=p��ݿ��rD 'G!`}���_ni3�R\B�'�g�4�;,^Ǚ�Z�r,s���՚���#�E�@�ߙ����x�#���	)��7��v�:�*�ٔ������? n�h��$�X��5;���plѪ�6�1��W���.�f[_�5�EXf�0R��Kִ�!1�`}x5����OU��Nf��=;�`߉�6��]%�Aޡ/�)��=�٤"D_v6TS��k�X��zw����G�u\0]P��h�C��O�ly󏅽��}0��6`����bK���&�F<�Ԭ��ݾ���I��b��m����ّ>bC<T�fW'I��-log�4����b��V�1�]�wj��M�{��ԭ��o�D��.' ٮ5��oa
5!��ɶa����r������(b��m��+:]D�m��?�9~�ʾ�?�`I�$��X�"����RX�M�8(�ZO~�Q�B{��K�U˅H����m����g��#�x<��4O�u��J�|G/�K4@'�(qm�h��<����l�Z�)��C�G�$:�ɬ�<��k�� *�'���l_�f7oG������J�{�)�}�0T���ơ2���}O]��h
�w{
�ԧ����VzI�b,�(�LAPvH$�'/�}��b!9ҧξ�ς�{��,toN���O�ekYl��y�Ƃڄ��B���]�B�]+�?���?�gɧ�Y�E��>�B��WE���٬K��`�8I!kЅ~��U ��ԭ��CkVN��%z�N)�-u��>D6Zßk�M�L��X&X F��yE#������ƻ�TAe��W�b�ٽ}~��9y��1x���5�H�(��9V���-�Po�f�6.�	��F��.�veJZ���Z�Y�q�7�ķ�w��
'���0�M"��:ݼ�Q�V~�����R��K�&{�:D��~D�N���u5�%���0�38�y����������!!�"�{���K�qmE�.�S1�76(���:�%������Q��#^�I�6!�a����p�g�qlT�T���T{5�Ҝt��Y�2�<)��R�Z۩��5�긍TG`ǳ��R��:{edG�c���G��ϗJ�g��'�J�^\�_@x��ɜ�3�F�T�K>�2;��b]��*�u��O3�Yt̢�s(U౛��q������9NOo������{u����EvfN(x�;����\6bP��*�>��S����̮9�Z`8��xSp���	No��$y�/V" �nkZ��d�����^sL �0��K*����h"�[��y`DJ���1��P��A_d�Sm��UO�j�M�
�>.G>foN���Yb����n�
�E���x����6C��EX�Uԑ��n���>��ap&��7��R4��`�tY���Lv���_,�8��N��Y��wϳ:��:N����������*�������}o;���SG�'��^cmu_)+BD�~��RY����㡡'��WYM��'/��FU`���,�����w̧�sI~(T�n`�ti�����/�g%ي�w5��Y�m�B���k�R���*}%3?���ĻlP�T���1hR�>��fʀ���z4��H����;�x�����eMu{1���u�c�ݨ0g[nA�E�O� �D=�r?���	�̛Di�2�X�������(>�
�m���Pv?<�������E帇ۥR�v�)O~�3�U���}��0�u�����B����ţ� V�����d}h�� ^ت�^�F��)
*RKFY�1�2[�C�ῆ���wa��t�i�jÃ��x���75�_�c9��식���f�8K�'��g��;�l���{��������y-�w�K5+�H����0c��;�pץ�q������^�*�e!_��H梂�'�"�+���Ј��SQԱ�Kaa�jW��`�����'9��ǈ�ˮ�D�7R���6�ʢ�V~z�Ǳ�������UHl��N���J�J���R\�r�'*��6iF	R �3����z_aX8���m͑F�踡��|�0|�a0��� �_/g�s��5��c�����姘.1�w����?�5�t�@�,�i������j4�[,�O��1v<(�浔p��?I �Uh&W��A�h�A]�_u��t�u��"���}�ǅ�K�WܙO���=�I�|)�ʝ�rC��6�#���q�@�K�S��#��T�U]���s�b V�'�0gۈC4i��	�@��x�8�~b����/(��1u�B�¿vX�ʶJ}FI�#��2�mF{|���:A|e)^�Uѯ���c��2�z�(d��Pc�:��Sˮ�83���Yc�bL_���ˡbT�6��Z��_������2��k�t
�rg�hv*��ʡ���]�<���A{Y�S�ì���%�d�ET�lIg�N�J�B (fY���gĵ=�{�`-�ٱ�B���قT�.��"���z+�]50�5�⮨ �z���U��%���&����p *��"��|��k� ��ޠ��F@R���� ��
�x�xڃ�7��ا`=��OV�jB�[*�q�1�>�+&��s0�������|�WVC�ـ�vu �)=�9�x�)wLR:ހxD|��	"��Pr�3�b��t��z��o+�6�>Ç���ӫE^m�H�w�?%/F��[����'G�ċ͚����vv����A� <�SHh9�c᳇�q��0E�)R�i�!iI)�}�B��;�����q�H���rD�~NfW��ݐ���
	�f���f� 3G�k���ZH�n��ٓ�Pp�'U�"�OkFߌJ6�n���I�C��������
E�� (2[�>ǀ��j��m���8�,��Õ���)�}��=�P�V�A�ʹ^E��P�S�R�w�ᝦ/m<PI��I�p5�#��R���G��uفJͯ��z��i�\�-G��@�-�;��UM���!�c�V�������b���Wx�g���,6-GSZd�4hK�r"�Q�:�$y�~�Sl0���а�-Nw�c��{�b�~���!�X�U��"勴bv����~=i���xs>��l���sD)q�$G6���׍I�F]0�?s�Jm��$a��g$f��@�V�+$=䪮7I�+M�2mnd<(`�Ɂ�� mŶXI��!_��K}aZ�i���W�*,4�}=��G�
i��cgf	 G͌�[S�� ���_��ѻ��P�93�~k�2n�J�?:��^���/f'�'ԭ���Ƀ�H��&������6t�:�/2�E�}P��3������S�cY(�j�`<�8s3먤^�5=�mk%�|���A�����(MZ1v�����Uk2�}E�ER��k3.�L��O�g�Ȅ���_��s�}������%�o�ż����Ճ��K�O#��V�������X��@E�H�VF�h�T�]6����C�^IsgE���n�[�&t^��{�bu���U���7:"��xi�e��,KE������\4O���H�KK��:�U
ǂ|�d=a�C{%&��}�<'M��.�v_bu�>4U�Bk�{�:�x��x�f 7�jk��S�Z�v�jb).Mj���ta��d�y��_�\�`�4U�0rcIֹ�E����#�>��57�{�0�M�xj���ISт��
��L�,��3vN�K����>�1�' s䟀�����rK?�{�h�x(�@�"`��_~V@5���zy_c�Uh���|�;��f������N���E ���ɟ�K~z~������Z2�K1TT9��ʷ.3S���@����Q�K���a�u��p�&��1�a�	2�և�Aڨr ./�����΃Z�
8�(�D��h�>;������5;+�>�f|��M�,弸 �Ȃ��|����4Nm�oHz����
	&�k�t���� �UV�(V�JkZl������}���a��f#��9Fʩ}@��^ED-سB���*&��W6��0I�Vgѥ�d}�|�B9�w�M�e�?T�� �-z̢�|CA#%rt�)��ŏh]>tUAc3�,�Ǒ>��!���F�Jn����1M�ШgS��>��TG`t�c�r���»�˄��zW���q��Ska�Z(zH���Y�w��;��V��������x��IW9_��3��1l��:@�ǧ�J��d�j��4iW�^Q�Cx.���\��HX7���|�� {�٪�o�������
��p�5�ű��	�{)�tH����2K`6�5���l���oE�T�񃣤��^o Ǽ�He��-��!���5���-w�[��z��M�~��{�h%����~�&�b?�UFu4������-�g�*�=�{)�������w�wK��<J�4d�`�}< �j�$#1�*��J-߁� P�*K�*yo�|��`S:��r^�X�Bؕ�=�:D_��h�Ľ�K-�&� ����eC�(U	�x��K�e�'9K��}:$�Ohc�^u�gӆ��~�Nq�%6�dd�e�8Y�F�,��w����[ϓD,�_Y =��F3Dh	_��t\̠@����]�Hi2�A|�M�>y2;�FC��)�%a:����� ��)Q���4�#a(�(it��Gq_|��Z�����Ͳ�Xfy3W��	R%5�~l�x�农w��ט��_b�_�ͫ�������7��'�T���~Ϡ��
�aŉ��d+�%���
T�@��p����e���f7$IU 'J�<[��RL_hE]���1�������m;� n�MW�|4�\�R��>7�p�S@�S=��Y�(mG����^�Bp W̢	�$w>�'-k�r��*�L�.�޲��@T�)��b!pܙ�����ĭ���7U��E� �v�ܧ����ݿ4o_a_2a!q�wL>))�Q����ut6��J�.���V�k�e�)��_�nh��66��25_Y�����o�N��MTP=�'N��r}U���Ѫ�%!�S}�:� �^DJ�-`��X�zy;�s��} 3N�wT�v{��~�m��a�#�W`Q�(�Z��*�� r��}��p�UP��������&���(�g{j�y?�H.�e`�Ȣ��{q��>����s�.�@���Go�1�Tt&~ȭ/1Y�8��`�����~D�jS�-g������N��KRV�e���4�k�M}���ـ�����6���93��7$o�}ڔ��
T#��<�M���p�	���^�`�w�E�IO�'�k�q���v�A�@�ZJ����GObܙ��xJL�=k�1/
�=gh�<[�/(�[��J�Y��v=�?�;����Xv��i��P|��j�U�l�G�i`����`4�2�oD��% �r�Z����,y�U ��Ni�o�FUFp����;!���Ye{�b,k��\�6T��c�3���lp�?g۬
�d�>�M���BݖJ#{���K���( �j��G�M���}��F5���#MJ�dր�d�'Ծ�U�X��J
���#�Gcd�Ϟ�xe.��B�3%^���{�Ϟ�<���b�9��摚�rbP\���~k���)̀(q�.Ƹ2��![�#��ߣ:��8�S��V|	����3l�dS�,"��6^%$ɮ!��7�Y!<4�V���˲�V�s�_Q��*���+`?�8����ni�.�,I��s4K9�X�Y�q���6�O�vt�a;A<����9ϔAv|Gm.�A��� ���ѨUiUHj�v�e�@�& %�v<��{0b�1�{]"+ݐ:f��)��������rͥY�8N	�>O�V@C����H�Ӡ��H�į��o�������]��uF�D����ܗ!`���u�! �jO�:y*]��s6����P5TT�����Ĕ"ٳ�t�5@�7	|�Y�]�k�W�����1�6�t�H��f�A�k2D��F����i�^�Q����T.�}}S��ޟf@C)%�:�nE�3KʉE���}&¿�q�a��.�>L�k����c�N4�p�C(3���� �OMh�ΧJ��j9G���y|�C����V/Q�
�c��#�;�d���t�s�@Rd�.f'"��4fO�=!!��`yP������[(�l"�U���$�6Q����kU�1O�ޔ%A�Ī��݌���d:j/ ����/f�ysG��#����S�����6�G��;���ç�A���p��fb�����Wk��%�]��'� ���j�`<���ף6��l�(d���S��-i�0��	cr��0����J�:�.���P��;�ɕQ�����3�# t/�mZ"��4���-��=�P��2�k���N<.:Wk9���rzZ!�Ï�i��4��j����WD���J�&�z[=g�|���ʡF cJ�����~J^��rb#��V��;!����T���8�m�	���U:t=�Q%5Qj��c�ڔ��~����!�&�
�u��;��B�%���炢o�{X�A���(�/��N��3��. 2:��tqq^ܒ����T��*��:�"�dt +ǯ�"�@I�:�i:C��F�Q��x�>o?���aK�'��H�̿��|Կn�h�+�EE��G�D�%�G?��m�'�����.S��(�t7���1�i/���w���D�7s�1������o9�c*u���Kv"���>�i؀�ȬN���^?�4�L|���z�K"ҦJ����.&��ʥ��C�s�����쀾�C�e�]�/9,y�E���`���Зh
\![��٨,�СB�'P��f6M.O��M��468��Ab�Z��P�8T�t<{i�.�C�ڗ����̈\ki�:������2@� t0�Q���|�"ߖec�|6G}P��9�����X�^׹m�_�=\��aQ=OK����C� �z0?�V�R�+�]j��&v�]�-S��-��b���Y���`�M��J����]{Wמ�/F,�[�+�s��D���U�����a��</����[[_G�pV���YyMd��A���8�J��c��ҴZ�2�tΚ��nYbĳhR/�$ cÆ
�;Lb��1]��Y�D���L�۸5. ��L��ZuM��=Q�@8LG~��W��p���s{�z�Q�\�DX�3�ʨ
�a�2מ�'HA�F�I?]t֦uo�}���G���~�������SX�3`@ԻW�i��	ԧ��}� �8���c͇�J�_]k��"���=���N|��8�AO%��hG�ֶPJwS@t,�R���D�8A�qD����L��'ayz������P��}��q�H#]��nm9�_�o���(n���ˤ�B}0�����KQ��ć.�ÑGɾ�p�V؋��05L�:���8���sԽA�R	�>sR}��r��w�$<�}A��F�0���ê.�<I����	�2rF�Yv�[5��]6؆��^�K��\�k���qy���@���q8�KK��g2�_hUj�c���[p��2�R���+���^h�j�[���Y_B�%�|95�7VqB�ȹ��]p-��9�O�=���)s0��������㏌��	_�wj����=����������-�U�Ȟ�����>����c�����-3�.��x� ��ƨn,�1T�2V�`�w�DR��ξ �x��:?�%g"kg7T�������\m�>gqs��y�(!g>��\���tUmG}!�nlMz�.̸J:�Z�%�K��U��: �%N���c`W���TeȒ}_�� <ؔ{�=;��b�>bそ�f(fHh����D����BdƏ�y��
,J ���
�\��@���HN��v�Y��$=��ZKQ֎�wz0
'gJ^�}�d-����r�<X��?u�,�����Es�	���~�����`-B���U@S���7^#*-@.�g�f6z:�)Kܟ�C+���x�vs�[��Ƅ�AB�-d���o�x?\�9�#�5�3�s�2Z�dk�rf��2&�-j���t6r�w�(�Z���!�vEG��ћU�0~K~�ls�8��vҦJ)�Q�?�<�4R`���c�������j*%��TC���싅 ��L)ǜ1�<�5�b��sb�1��PY�Mp�b��!_�������}�?m�����0���Z@�F�\b����q�V�s��V�I��S���a�B&���@+�yj�W����9�����=�y!.&���W�C5i#������� ?Vpz�~r���Y��ʶ������Df���
B���{�t�4V$�
�����B>;��[<#�$��r��̭�ͻ��~��m�}t.�$4�vU�����;s���t�߳[K��Y>�-z*D=H;�2���!?���d;�����a�q˵�]J�s��_*�4��O��_d!���䔨<�[!�)Ŋ�h���L�'慠���aU3R�p�uB @@����� �܁BO�������#$dR9��¡�7�5H�
�Z�0yx��1F�.g�"�@�\��o;(3��؟}�E�:!s��DSy�V�R����ϸ&�Ղ?�}}CϹS
J~ץ�+������;�: v���%yYj�J��v�8�oy}���F���N��&�bͬ�5>����������}�<��T����D��=��C�e�6������ֲ[��֌o�o�h��	.?�Ί|�z�jO�d�����~aW/ � 
3�z(��O��{3Y�xy�|�;l���X�p_�v�0f�kK/�/���x� ~>;DkVh	X���N0K��>�6[ހؗ"�3֤R � T��ƬȦ�����k왢�K�����:H��R�x�8��B�ԏU�@�}�	�;����ɓ�]���p����?_`�0fB�/J�4�<#�_���W���t����%	%4+T:�7�e5�f��7!�mpu�Z����m��_צ;�`�I��� �Զ����a���n�B�����W���.���,��g�o`.�Ԯ�@uL�)��K�z�W˷�k�����axf����Bi� ����-_N��K�{�EB�y�����JkS#�%~�k�����S �k-����&h?BuN��W?Hl<����
�R0A�����	�%�n]���vRT��01���������\�cp@�7{������KU���Jd�3c����!�Gȫ��V�|�mD�ND����m�)V��K���hH| �g��.�=������fؼ��CTX$d�z���62��|
����9�)�d
8��\�.̟�������Y��Y�mj����T�ҥ��8�w�Zq�F��� �G�f�/X(y���S��/?��L�E.X:Wٸܩ��[<�{{"��mK�h�*��/߆�J?�L�y�qč%�3�\^�7(tdA����@��J�;�F�9��Iش���AL�mZ�(�O�)X=˘�~�)�{���|=��΀��fStU͒��}E7�-��x\u�r�R�8�z{[M��-C����z7,�}ْ�D�v4.�Xʏ�Nc�+)�ػ�CKK�\y�^Nޫ�p`&W�oO}>�)�hzR᪓����	�I̶���!�ݩ`�绯#Zt��o0y�zFS��>Щ��$������X��#ڭ�?��{��bI����"Ń,���هm���^��Vb�O���_>����3, ?��y�C�f�E��U��$��܁\��q\ǎ�֠�f��[�ſ�m�Hs�o@��8�k>��+ ,�IO3�o"��E�~-Q�u����@�]?�__)K~E�Fe����os:���Q4�t���"�+!��
JR�Bķ�a܇5��@](�k�O���:�n���M�ye(![��!�9QK���H��N��z����	,Lh6(�w}�;�Q�Uޅj�PL�OGD����'�!�+��%�
ͥ���)O֩�k����o�T��n�T��I����FB;-�d�b4�w�*iU��u��x��@�jeK����@��l� Ȗ1�����#9#'�G����۠��ص��8�>4W"�M����j����샎�{���6&S׫�SXϨ��ߖZb����G��A{*�i�:�C<����:��yS�bw;�q\,j\4�6h�c�$��Iv�]{Li���M���집��bP���-����`�84¼\RB��x6�h��$q�g� �i���!����H����!w� ��bU�OX��1協���Y�$"#�����s�6'e�u�L��u�'�>`VRmq�Q|�hnU㰬����u�]"j|t<��`F.K�;�-3T^�̃V�VY���C]O>�ȡ)�m�#���IŒ_�@�nmY[3�t3�	�,�� ����m >�*�tv��X	���PI�N^�c�f)�+a�A�����<�ǺD����#1�r��t�&=}����e'��NϿ��I�5��8ЗٰL�<Mô��	���k�!C<�-3Cv��S�`c�Ez�@�_�b�������nCI��陮LL��E�9��1��i���C�E�M����/��a�ĝ���g$`]�k��>���)�����������[K�8j](�a����M,9�@�"2.����X~����/���
l��v�_�I�����e���ݼ�������H֝��0�V���oV9��q�{[�v�����"+eY�?�CZK&IM���q�����s�Ao��t�8����$(�#���;`���KS�;����O5\�詿G<�o�ܱh0��w�M��z�c얔%�$�`�2�'��KP��67�����\xZ���K���x����!S� ��<VO��zE��M%K�AX#S�>O0{�u�A�Jp��C��U�L��H#�*j�ha�<�^�+H��~@��؉m��=�/�SJ�>�/p���~E����Z�L�|i�rS�������
�, �X;+�7�y߄N��_�WU�hҹr:.��;?虸�D�T	�= ʊm��l�_���5C^��a������+'����m��/�y��-�ne0?���8���'�YM���h�0�6h����O��8����;� ~�G��Ƚ�;��H�i�}�:�4[������Mv��&�k�7ȣ(�/����/��1S�*�SB�q�O�s�u�>@�L��9��Tw���^v!�N�ʮ[�H������mE}[sj�xCV�2�^�k�G�`i�Ng!mv�'��ke���Vl��$�C�2`���L���F!?fiQW� �|Žx�V�7�M�}�2�?�hE,v=�L8's�1�����ʉ5L��n�f���"����<UFc_�țK�Ƹ�������ñ�)�1�*0ˬ�8�d�b����9mgI�`��7�{tj�y��w��x��K��RZn���j��p�pR{�M6>xu�7��|j�>���)2Y�/<k�M�&�C�Aj��a}97�~����t� ����yyn[-�;i� O��z-!�.���)�ƸA�Ag�X����no%����H�X� �**����֯O�bAPݩ���>�����_(?��XjX*����=�;�e�bW�j��kA�~Z�K#�ٵH�;����_�e��㖴Z$� �H�+.�c~kE�m�Mh��$���B�@* �wYM�E�w���"W��>�O���lji$�-{�4�Q����Z6�HCp���
~��^�ɲV.�ʲ[qqN}�/�pF�݌��dɰG�=� ��x���������J��V�8i�=�'$+JL[O���9CӨ�Ƈ���C�I�*e�Iۇ:�z�f�~(���	AA����G��P�M�MӞ�g6����kd3��,�4f�w̓�&S*���hœ�{I��fe%�i�EE�)މ�Tv6`6�h��5�iЪ2n6�b���M��2�F�k���J�_��'UB�\G����M��RR�Ҍ�+�0Ίn"��M�0b���#�&�\<�
������I�"f��$�W2� O������b_��%�RzD.�ٲk��|�[�]&���>+��hΘvz��ɇM�rh��gh� �ő^���W����r�`�QE��G�E���~I�ᢅ�.�H��z� k�u�4�Lt�����>g��9Z3�i�]�M�6,���)I?a�,����:�������������w ��2��5�d�ͪ���E:���
.�+cЪ4/̡q
�0���9���"�����js��Ħ������G�QA.#��n띘�&R��!�p��������a��8��|��3�a�u������CUx��Y�i�R��UbqT�Q�����D�j�.gNI3�ަ��<���WiǞ #�ͽ���;��ؖ����m!~��`C�DKq��7�pֆ-���>o�A=�_�]��j8K�<hP�%pS����D������7�� ><`�|y�1�����g06ZmZ�tK�Q7���G���Xdc�O�v�����u~�G��7�H4��|`���v�I��<V[�*��Σ�|�t��w!H�ʰw��N7u�[�1��O���=�#�J�y�{��"�K�ŷ�j�a Td��
p~X��.�;�wB=@�U����g�R�ly�'V�,fXø�.�p�
��~��=D飰�G�F�nG� `�o�C �x33���(��MԹRV X7����i"WJόZ�{~�Ӕ��0p�&m�ͭ}��f���T!�^�� ��o'3d4"�]�iU���ΐx��{���"���]���N<��Z�:Ld`�u��O����I�G8֪�����y�j���F)DH�>��m�C�wѦ.����b-�7�ΌrX��TV���I���q�;�A }��:����h�F�<�IY3<1�ZH���n�v��\`:�w&%�1i��6�bTz��t�lS�nS���M���zB0���/�#(R������0ӂ���v��,���'�.R1�Tj��W]b�Mp>�/�Y�9-1sr;��&}H��[��_����ߏ�o�{�2;t���)��X ,�Q�K�їk���H�C��=�ņ��[ ��/w���|-�s���O��LA�p�1��~`BL�X)�]7R�����" aXz8��fQ��I|w�����0UB;X\{��s��~�[�b �^��<:m$����.�ͷC�����0�#�\j�B��϶��u��f���yZq+��w�X�O���	��> ���D8-AF���{�D%6�I��n��W�]\�U3H��xD���1��,w�gүΕ�5Ee���?�l� �xo݄s�g�����]j����5i����k����@��ˆ�i]~���]O{S���!��E0Nz��[Ts��!�s���̦'�~�Ɲ<
�����2mp�%�{�P�Y��:N�탠fv&,k��~M�͉����g3�*�����	�#R��ջ	�y\�����V��|�W#�E��K\�!gc��q}|��Ȥ���.P�8k ��%��؂#�U�|�I�O2�z���(����whP
���e�I҈�eՎ,� ��êXŊ��J1-�5����Xz|L�����pYF��mн�L\��2���*��*�HJ�(8���!;�\`���OWU L�vBtN�*5Ǳ r��~���9��ɑU#&@�U��n�[�#\Q��5�=���p$�!b8t4�5�I<y��c0< D]�,����!9-����n�Zla�,�6��o8��T"�o�,Uل����핫�/}f��q�����Z5�`�QY�B_�dntr�Nm�yi\P�e�8:0�(d�K���OD��Xõ�J~z��l��,���@N�o��B�kJC�6D� /�����}6���I�z��"��nJL�J�J&��Y��|��C��V����i��퀥����"�0�F���H�� ߛ���
��ٌ��r�
���Uo/�Sj�D��j�ڏ����ʵ�_h	.�e����tuc�W�1��[797"Q�i�\��zg�L�Ѥc�PemCм+H���|J��n�	�'��:�MR���=����u��S6jԹv^x�V���9-������T�B�F}	5�8ivt���V�&��?��$t,R��������k�)�Y
վaJ��n��ҹ����
����BYa�_BD�	_Iu�m͙�&� - -���)C��.�tM�62�g:���RǡX9@�Cք��� x�i��Șe�b �G��:JG��s�i�qJY�6��d�S�g$��}� *�3g��yJ�R��h��|԰��=��>���'�i !�ؖn�8�Dzޯ�p/D�y䊳�K�T_��a��@���}�#�o�Pj4��I欝nn���n�<��TG@�R�O���|e����+|]W�H�x	!��Q��0�{�����t�!�sc�k���\�ￕ�K���{�FT�?Xh��d�1�iW魽�y�Z��P�6�-�D�e� X˰
���.�{��|0#	UZ�R����R.}qܡ�|�I����~��Y#Xh�) ��ȭG��Vpza/�r������gHW���L��i�5_�-���Y��Զ��7����_�;�Qf|��)�5ă� b�of<$���{�)C%� z�`�墨!���7��k��	-L�
�
[!�?����
�[g>�Cɦ��!�k�]�mP��{z2��O�d����%��X)�D~������e�n�,��J>W^��^���">jy䫝�����j�ջ�@��V�&�+ي
�����5Xmo����vs�-o\�_Y;Wj��{��<�U���)r����ȱ�C���A�����⩨��o��^���יi�ŏ	�������:�u���j�r�[���;�y#���(����0��gu؅��VK�X�������W{I������ę��Gx<@�8���l4oqXD�rZ@4��%�92����#D	�s[�Qqï�yw{��e`�J�Q�H��Sqq=q�����������u�iN'��%G��
ɏ����虳Ns	�@5��������5;�5���T�O�b�^b��.��*����/�P����
��,���~�l6�ת�������,�oԈ�4�>xn����M�Iq�*�&� U�Jˉ%��oYޚ�S�}�͋�p������mk췸�OC��Z�է�a���0/�`�og�Ui-h�뇹M��=��F��!W�~����l����Sc]��?<ҳa���|�A�Q5���tvHG�G�֕tq���L�JJצ��S���RF�l+T�N +�% 2�� �^���n�|{P7v��'��@Tj2�*=\��~Z�w-�RCs�k1P�2�v��f��;���^ۑN@�I��T�z6H�=������J*�z�e�k�^��M|k�_�t�j5ZO,��G�r]Iѵ#ԥ@�6&5䙔���̙=���4�4^��T2�p��ٓg޴��-O�7ca��N�����u����)�F�܇�� �o\F}���t�*��`�<���U��o��uNsT��.fY��:_�
�F�ϹTT��@��M������M:�,:sG�6���@:���С���/�	E�`�X��A-|�+	,��[Lٺ�+g��Gi>zj�y�n����?����3+c	϶�(����D�H�>��l];��ܼ?�z���HV7PM_��w�i��<a�����CW1�#�ۋ��>a��t$���upC <�G�Iہ�a4s�B�S����.gC�8�� ��Ҽ��i�L:OX�S����μ��Xp�Q	�Z�7Yz� ����`Rfe�P���!�+"O�>�F%����i��9�(�f�cc�kOcD-���-8	�E$/�w���S��tf4�����_m�e�A�#�1�M@���ڤ&����t��źeQ�կoq���$�6����� �Զʜ2�P�9�������r�b��ia-�r�f9�^��S��FQ�����?�e	��@n3��͐��H����Q��H.O����&��� l�g~�&��������� ?4	b���g�0��"�ɧly�}ȟx>�7�)c��p���$��J��PU I���>��x���]�4���}�WL �6$灮�����~k�{2�.P`��앖���7���}�$ډ�U��k*���[_J�:�v3���H	��Sg�G�����❢�:�k*C0�I#�$��ȩ�Ɨfu���e��1w���A�ެ����Ze��E��d����_�FM�@n'�Pyp�Fa(�`����W\2���͒�ŨZ&���������:�(�-u���hH~*�o�h�����a`�s������`_��I�ͱj
��*�R��*���O��N{�K�%�ޟ#\g��Mh*S�Ӹ���Ϟ�/sCii�B��r�ҏP��a�]��1A��3AC��q@6ap���.��Tb�J2Q�"�������K@O�ogm�v����I���6Gz�l���'��iR��s�K�C�A�č���?O� K����51棸S���t>7z^�o�31&�tK13���e�]X��~NJx5�B�-v�7u�\IZh�o��Rб��"x�{c.��@��t� ��oA4���Qܬ,�w�Y/[&����jƑS��U��6:c�zez�q�r
��U��Hc���*�[־�w��/Q��v�.�BשL�۽����e!��&�ö.X�T��M|�@KTB�ݱpji�U8P`qߜ���QX�H��`..v�C� B'�a�����ˉ&���J�x�\��!Q��F�>j^�`T~��ݕ�G[��!oh�����I��0tt>1cO���R�����zЊ�U�7^Zr�|���:%�l��?���Y��m��^�F���[ܘ�MI���\?�:�Sغ�ͻ�:f�=�2����f�q.Pə �0��{ܶ�۠d��N�'ԖXa}��ǌ�΋�$:�z#F�}X%,N{D�8!�#�'%7��E,H
Q|���V%*H;��NB	�A�I@�	��g
�1�9P��s�-�rHT�2b[��&.����/4�I{���K6BU1a9nVӍ��f�ɨ
V�ɧ�"/g-���,xcn�Lx�3.��a�+R����N`���WcUx��\����Ul|w���� �N�ʈ:�J9��}��<�ݾY#��xM�A��`!xk��������;\kw��&��H$ᙎQ�K;��_52!k?�2d{Z˫Բ�����J��~����r��h)	�|ܦ�b"^e�8�%}̈����1I۠C߯��𤻇翜l�c��
�O��np#��9E��X ��D��'�.ǵ_C��b��i�m@����m������6��������Z�OcfY,T��
�p��J�?H�����.f����Ra��NCcҦLx��P������;a�'�C��t|jG��ׅ��A_���9g��w�!o�����z̋ϴyw����ќ��
dyx�p)�,6���kYs�.�D���q�1�F/��-����6gn���())`9S�1���鼪�&��������Qc{%x�,W]ފp����˹���2~��.օ6e��r=�̺�0җ�G�k��N�d鞨$Y~l�� �r%���� ��@77�d\���gLk�V��v�~�P�(�A=d�'p�Cܞ��Z�$)����ɤ��z?jן���5����Y �h�W
^`�DN�}`��x�$fQ��狀I���S`g��<E�mZAB�ޓ[�q�t(�pؑ��T��1u3L�%�e���,<t�,_@n)q�[Z�d�$�)W ���qT�f�xٰ��֘��.V�[v;kטY8��t�Vn��0s-E�M?n�S���ͩv{\N�&FhY�3~2𓬤�>�7�SP�^@T?3�e�/O桴^(�Or�F�yX�=$x��$�#���8 C�jyΦ(�k��n����!ف�\$����,�����Q92��å(���,ڴ
����h�"Z�c}���vbg��<j��wk�{��&P�g6���ء�sgK�.��4�i��u�Y
~̛o�p��>�J7�J��
��F�Jא05�%��G�៉ή��,	���i4n���Y��$v�����������(c}~�5Ƶ�$s|l��Yj�x��_opg�ɮ첗۵�˼�I��e�V����9ԛn[�{�~�W�L�L&��v<��W���q���o)�[#������ⲛੲ��\��l�G�YB?ٺ�p
Y��}'�A�E�9��u��ş�&G�/C��N#��u����J\<bj�MU?W�'���k��Ì�gm��d)Oqat:5�Z>طa���8��ɞ���OD����]{�4Պ+ǿ��.�#f���n*�F�{�sj����)�8p3�O[q/NH�yqJq�:�������2��>K��c�����b�Bh|{�vd<$տ~,w��2E�OI1�+k����i돹�Cl��\���zD��0ctp~�q^ү&����乭)�����|h�o΢~_��M�*�3��uU�F8�
$�9eߋ��c�E_#���F19^�ӥ�BN���q� sGF:D����O�E���O~2묑�֦4w¤F������تB�VRˏJ�����1A[���٤̏�wf��V;��f�ǣ!�>�f��b�b�&���6�{������K��j̢h�P�="�w3`fd��- �Z� uv>��#�r�����D�~��r�M�2%&q��L'74h�kHU��|��z��3M������"ͨ��.�����OlDW{d3�W��_��}
�v=�$��"�DNr�#��p�x����9���������%s��48�_B�=��H����Z��6�����1�
�,V|r�S�V�2��X<ܿ[�K�蟖ݒL<Ά����I��L��<�5���%�t�'�௃�3y��$y��;�Ky7�I�(�M��m�d^�~�@CB�ͬc��Q(+��2~�bNV��tB%{����]�t�4���P[x�&m�Z�d��i�C]1�rX���q�K^N�.��Tz'�\�B�m���SoE�
ڣ�q*�:�H���-�h{�HU�}�(5C3�)�Ϋta�̅t�ɳ�]M)6��~�J��G��f���p�՜��	�{�(����v�J94�g��.�&a�����#���ԑ�Vq����;���<�9L���������:X$癄���=�'A�dkcS�L�ʗ�0lP��R�i�:]��,�g=�����у�?д�@8��k|��
�І�x��:�i$�ߝX����.���S�� �_P�0��%��Rh�np�7���oP��$Y�&#iӹ	������hT��aь��9j�)i�)����n����֮�or��r�1�I�n>�)��;�x��*��r�I���l�E9�̽��_F�6v�TX\���~�C�r��6���	q���.�?���'�R���U,?^�pv�)R�C��Y�r�&����;�nr�α�f�W�I5٤��<އ^���x�p2y����5��)�Q�K�eF����rbp��U`ite� ��^��`��E6 �8_W�� b4���┺s��t���cF�A���=\�h�F�����`Y�"cH-�9 ��{6��Z:H9Z���8#����3�c����?nDCt��)��%S�$���q0q���Szᄵ�ަ�@��M��ߨ��`{�D���9�v3~;.e�g���/˕s��������*��ƅ=a��͏�FsG��9��eښ ���-�-J�n8푞���z���umH�[�~$��%��`+]u.i^r/~�\��F��y��?@L�9���:��Eπ3�&`��!^��V� �K�m�����0�*k����l0��3��ڒx��њ��b�9��Ud��x������!���z�2Y��v�Ŷ{êT�O�8l�����S\q:�� ;�KU��9���5Y��]JNCe�/����UH�8�3��Y��I�x�-�ξ(hlǺ�Pσ�5
��4�I�l�X~������±aT��-�tQ@ѹL�2�"/p����7�$��:�����H:�(�a�ʅ2z�'�=�O<q���0�Hb<���-���)̵��,�31f� �S4��0Ιa�`&or���L��Lh60���@3��h���Y�v�� ���k��X��{�A4��E�@� ��o5m�SAr��lۮ�F��
�R���b�6?����ѫ�':�B���7l���?O�.�V��j���x�EO�#�9y�5b��������ՋnP�����9z�^//l��ڕ��������&��GZoT��l.p�h�-�!��$�������~A�i�Q���M"��<�<J� ���ScVQ�ɳ��C����md�0"
u�3������z�N�Ӷv����N'8\��1��� ��*෰�r���n�Љw{qX�$G��n�,C�H�:����S24\�P
+��R��*��m��W�87޳�ǥŭ�ǁ�}�S R0����-����3�t9"}�-��&�M(���� ��qs"�dȄ���~d[����Eo%�ȋ��o�E� �g%�A���s�*i���ֵ�׎9��_Z�&Ƣ����-$�*d�@���ֳ:z�_��7�k�2=E�� ӆ�|p��U��[�|�Q�~Fj [�X�w۝�OA%����5�ć-�s��2����3bcN����q��K�>B��Z'Y[�q�L��`�ծ���⭇�Ͷnr/;���P@��-o�X�Cc����n�+l4����LH��楥�{��w�g����t����&H�N�܏P���\�J��ᮑN7i���:<��wf-�"I`�<��\v��+٭I�$�i�}泠(�%l�bY�~��M�W�LE����>�PI?F~S�������EU�%ΰ��l��S�A�Q7��mt�=�AV8 j1�!}��7�l9���_��jp��5��d@����1в;���Gַd�~��\E<�bm�Ӑ�4�����%g���-��kY@�MRS(t�Ks���4�Q��~��#�	��;�R���1X|�7ڑ���$�ga<RU�L4��!,��OK?��ώ)�T"��i���nIS@��s�3x<k1O|(���tI�˝���r{ۧ�]zr�^F2.�#CbP�h/�?��P�:"i�%oLã�u�����g@�[����l�n<�ϸGAAp�Z�u��{N��Y�ƕ��m�.�߾f<�����e~#xg�`3Z؜���5�X��B�^Y�A�t^e�x�B�)OA8�ݔc�]Iծ�e7�^%�4{6xX8>Ѡ]�U��TG��!V�B ���'�ں��6&M��BI��'j3�R@���!j��,�$0T����Xs�C����z�<�;f�Jyblٱ#A�����d���ȗ���m�>,)�iPæ��B�%l=�w�{_�����L'�Ga��|�l��!=��� ��u��r��	����ˆ��*z�=M�W�,�u�(`JC��b��O�.(�J��pn��w�kV�T�,�r[���M� m��i� C�΋x���P����lH�Aѽ �tJ��c3����e���C萰��^�E�"4���!�&�ҧ�vL.���"���K�?	���@f�>�o"�1�m�֊*o�c��`�RQ%Y��1��ϵi�%����r�b�ץ��*�����������˲V�Լ�V��"��7�8lK���DP���ƈ��_��-���b&a���|N�k�4+�CjX��T�Ox"Ո�f��R�M�q�;+��K�ԼԚ����]A[&�jFŌ5̍��IsN4��^|
�޴�d�6�7 �K$����HԿ�]D��A������)*�-s�H�*D�(�ʇ�h5��8��(�߸���Lm�z�J{��sX���$t�͒�����knw���󵈚�6}8k���<y|Rz�{MŊ!�܃��p3ʼ�tL����?�Xm�������)%Ǥ[�X9�bRB�!�~3�]�/^��O4}�c����V�Γ���SFeo��-��S�o��0Pzp�����B�ŦNjTdgK=��G�b�v��e�e=COIv	;�0��@!���b�]������V7�7�
|_���Uih�z=5?���|����֡G�g3�Q4��"���{��^�A����*P�,��{�ύ~�.�O�>�)ʍK��֤P�[Cv����%k�Vj����`��줮����a �8wnt�N�j��̻E���b���j>Je���{B)�����/L�����%�/����税�[����i,;���f�w%�uu}��H���ŉ�l!�E�~��.â��и
1��#Й�g�p"���Ѹ|��w�M�xd�YR]RpU�buL�{��~
��"��O�;�b+�)q�D ���+U��t�L0��Ɲ���6��O�#�jc���ꔿ�����ؒ�q�0mȄ�xh��>I<�6өw(e�%�x��d��5��Ί��ףʬ�a|1���#� ����S��;3��:��_d����DQ6��G����Y�X a�ƃx �$&0�0p�l��ܱ����������//3�"4�EUnLӪSP�V=/>���u�R�:��;Z�e��m,�D�mS�6���$G��a"�oB����D7�ctw�m�i 
=t���޸��`
�(fЬQ�{�z�\���D:f�m]U�`QDi'Wr�N�L*R٤�]IUa�,F{7�V�{�Ck�Vq���Y~����7���Hz�T��6��J4aJN��rL�B�p�p/���L�VT�1�0��0��v��^��K؎k]��:�	j��É��X/�=���XK�'��@�&���"殺�5��{Ɂ�zbh(>Vε�TKf�79���^�Ǻ�y*�������;y�塹�άR�}G�KT���"�G�P�ŲYk��Q����;�8A+ZLY��/v_�����g�ᝣ�_�4���}w#�^�O���N�gv���Ô��N��+�B �Vn�`{�6�H� (-���Ff�tg ۹�ڕi�`W�ߏ��q����|t���K��fVΥj@�/�����\a1���ܵ;������.�&\����J4�a��V�cO�,4vImw�;�i�TՂ�>��i���:����)h�Y��'���r��Po�6�h>JI����+ʩ��V9no��L��8`m}V��KĨ�TU�Vs���3�cR���cDԕ�4�Z�:�
��F�7�}��KiV���'���]���H��D�W������M��E�{$@�)�I)988IW�/v@4}X��9��B@��-*[���/滛�	Q�ֿb�M��m����Co��W�ɞm5O/�7�:₲%b�G�y gF�+t�3�QӉ��ʪ����/�(�9�yub?�b��s5��W���s��N�'��-�����|$E^)Z��E<�:����Z��
xwh!�9N�PA}�Sy/�������hآ�6ޝZn_�j���g�i3˗H2��ڋܬs�k��P��:a�����=�m��| Z`5���h�t��W#b7?	�d`}Cp��X�������dS}����&�$��J�k$��F�>��Ud5�~l�(����19;$��.�f���:�.��5�-�����V�ǅ0c�~� ������6��'8�V���q\�"� ߥ�{
pL�D���&Q^{|]�-#9�/Y�(�^��B>��M[�c3A��T"���z��:)B�<vN5�x��.���-��H�_��|�(��b�"�a������:E�
�헔K$,òŘ��d���5q��VC\0���Ϛ!c��C�?D4O��C8���i6����r�Щ'gX�+��C������)-<r���������#��w�r�S~��젷u�ޑy�ѩ�ZL#�j���e���Ԩ�����L|N�ҭ}��s��j��֐����w�G�pa�c?�8/Ĉ�H��͇�M������!��-��']�E4Ԯ�P�ie�p��%�s�m�}��;'O�&�M/2'J�R��w���C.5+����6���X�1`f��@��j3�M|(�*]߅%{�X�RY'J��+�O�yp�]�G+t��v��[�0s3"Ƙ��4��e[\D��j���_q���N�֏,�����5��S�L��ſةm+�s,��|@e�Mc(N�7�[�z�U��R�O�bٮd´�6��4T
��������GZ��B�GZ����@D����s}1l�����9�� �-p����wa~�<P��!��3V�ǀ/H3t�Ց�lw��N�i���hs��5f�k�����ߢc��������KNƽ�dʫ`�%�Y��:�6��	�5XNJ�u6N<�a�2G#z��{��㳎#`���p>�+�e���ِR@�ƈӽ��%`�#=��sJ�(E��j��]�x!�<tC��9	�i�j��0�k�*������Z�|���3�EߓI"������B�����h8}N�a�K�k���G@�� 8W�U
�2jv��#�P~w�b^K������ч��,��O#譋#!��y�L��Op�4&���B�BZb�O����r�-�=i���[��Ӵ������A��P�#�~��};��2Ґw��S!K{��� ɋw��mӘ�63�DL����r��i�@v��i����»�ۋ���V�ղ?���vy��s�i�yAb$F�Nt
XP��h�1X��-�M	�"�E��~�&����M���f3�FB���N��W3㠻���EM-�S�C��iz0�B�H@Ǔ�{��!yں~��>�f{�Q��r�����ac������i�����s5�vEA�O�h]5���m�$�+�
��4#y���S|W�+����s��&��#�=��y���p��B���dO��������8���Y*	#1����{�]dGLM�6δ���G�ቴb�bϝ1g�u�v�X�h�a.��WؑVK�;gx�b�4��+c#Xa[WI5L}�ݮ"A�ox�ȎN��G
~x�����#��zF/F$��.jxE�O�����T�U����V��0�({�!��ܽ��]0�����3��=�Ő\RND�k�B[&4��܅��P�7R��]b�舫��=O���Z�b��6﶑��7X b���ݛ1�ݕC�"��	��l���? JX��_�e���8^4v�J}��L\�7�Z��Vp�8 yk=�E^e�cӎ<�葨�`�L���3���f�9s<��H��\<�Y�ҺHp���;��/~c��p�5m��:c9�N\4�9�z�:����N3�$���8tտf9~�R�傿��v���I��J�W�5��c=�ʃ��خfL��$�|7�?��l�J������~M&�Ŀ����8�`sP}����i�W)���Aˇ���-�<�8?�27jμۓȦ�����v�:��ⲉ��J����֐��z]hb��gSd@N��J��ۜ�N�h;lq\X����?�l� _u���[��O����,���u�X�V��Q��Sᮌ�7��m �F�Q�\��ȗ�p��y*���~B�1�2vxB�\AG�ѻ�zs�ù���Z�}s�i��FZ����ٶ�(_[��g�r����`�>,�.�[Q��&H�����&�;��.A��FZ�[� �ʮ.��&v��FNM�F�r���f���/.!'u��吻1Dq� j�v�Y�9�A!a�´F�D�3?�2�)�4��~@ҙ��w.�����6���_���c�?C��(�3�Ɣ�Ԍi��rG�`d�~��z�
�ڱ���|S����5��Ӓ&1�o��K��B�-�?���ަ�X��rZ|{��[�� ��.�ό�`���6��̓�5��;�[���7���N�����T`F>�f���~i����z��8���4�'��Rt��RƎN��������̏����7�dŰ�o�z�sLwe��I�)�F��N�_قUO�l��9�pz@�����q�r��������q�u~���m����,�� ������Lw���-q��۳PuK���<�DOǫ�%�Hw7h�v�z�?�V�懓+#��{m`:��+C�%VI�nG����y�"9�A����US��~��Zk��8I��zߦ�M\���/��A�[,�I!d�翘L�>�n��TqƉ5,�k��,�����^����=P��qq��U�EՐ�f|��y�3�yT�hX���^��Tl��-�c���@����Gv���?%ꘗm�)U��/�H���epYJNdG�bB���/�5��"y�g�岴��
"�v�����*c����@㭋�Lc�ֳ�:7��2���E��kV����a��1�Kܶ�UĴ�
 S?6���ƒ�gB��מ�T��joh�����c�@ǗZTL��mSF���<*�b^�z�7\"v���`�TWJ7���o��x�
m�Q��윿�9Q}���g�	��z���Y%�`1����U��$����X �0L#r�XV
��B'hq�pCFA�_ug7��';U\��/�<X�=o�w�c��D5�u���;���[��ȸA��2�K� �RM�z���U��J}�*[���;㌷+d{aL��C@H��N��p��g���ka��IK��0��܂1�=���͆Kqr,_5�$,���Q����ە]!/T)���D��'���PH�B%�5r�x+M�H��9�bfP+�Ǳ�O��]�RL:c)^� ���c�|U�z�F�"�縮+@��fY���{�Z aU�����5��Yw�I7xV�v(ޓ��c�LJ�L1Sai`o�����4��	��}.@�K��	�|[�lP��Z�^��K��W0�P90���Q�ߝ���}8�������j������TnJL	�3�ǈ|�k6U�8��.o83n�>3�5�'����ܐ��t�)	7��l[��*�Ν�[��tl"q#���"�˦N��R�Q�[�w+63s�a�b�;��RÌ.�z���m3EE�<�¬�4K$
�|�j���"x�Mx�7~�e�يQ�/����5Vv����F�\8�&o��s[���t��S���y����A���=�TA{��ߖ����W��V
��k%(�U���z����Bi@���ɠ�d/�*���G�c���Б��s�����E̟y�	�.PBoi+���%9rY�Fu��-���2��n���J� P��N��c#~����#�t%۪E$������XU���k�OZ�����J��zF�gd[�A�s(�T�wI�O�7N���-��~D�2�o�����%��c�����Qm�@��z��i�F2�	݆��o�=bO�I����9����%��Uk��~��l��I<���4XKE����\��(��L0�Z�s�P�,��4��lL�:8K�$� �I��t����q�E���S��=�C�5H��tLG
~+�YDE�gǾL��ys[�'����cl��^�ܙE���,>ً��E]-�����l������VG#��d�xJ����o�pd.�� �~�(\��]M�%��`��6G��em�r��qT���W��'"�lR{u��jm���%�Bui�Y:ٮ���@OT�{����"�t#�rpӢO�Oeu�oz+�@�|�)��bI��38���3ž>��Vu�W�����OѤx���� ���-5���-�>7㇜�D[wĻQHL�ϴ��7"�5�d	����в�)R�`P�nb�$���H�\%\�T6��ԕ*�F��M����3h-7p���ċ���7���Y2���@%&�#a�r}گe6�����\.b��>�;�X�*s�k҂��m�]�Y���UJ/B���Э�"�K�#ܤ��Bx��.ߛ�{uWT�]�?���K��՘��Ե�vL
N�!���+��Aұ���Hp6'^)8
�~Am�f<,�^�~*Up�s��8"�V���a�wzŰV=ma�ʱ�鏞�.�'(�s���Jk��S�c�D6p}�ڂ�z:�@n#j)��c �O��Adf�pF�*X��z���$�'c.jQt�e�[�<��;�j�%0z�k�U8VB���iO���/^?�}�=� n�|���Y��wq�}��ݗ���Mlk��39�⠲�U:4I�ٲW����g�tQ�8#�F�~�?�� ��~w���������JfB�";�z�Y�i��h�HJ��Z�����b�ٓ/��i]�����i��x�Y����l��\oj<RD*���ֆ��3L�y�T�����3�z������d?0�����`7�[���.\3���: ���Trܘ�K�
�4v�ɥT�ˡ-Z�ƭ�=�l$�,����Z�z��o�^��|�%It��w$�E�d_�8io���|���a�F��WWJ]���e+��A{=��;�@�g����~ m�Ŝ��.�B*�g��	�]�!����J�()l�`��h�p'ZDPC�R����W�\���n-��
�T낷��ӏ�*S�d�G0 �_���.�9���	��#I{y�X$xP�6���)�͒)8�e{���H]Q����}<K��G* �CwNF��Md��kc"���1��@Û��qw�rC"w��R�0�-�k-��Q��o ���?�t���������
k�������6��o�*�֍���'�7�3���,��D쬊 g���*�|W��O���d��w��M�0�ؗ7�3b(O��$��v�5X�{F�^k#�ٱ�YŁ7t�#X�D�nnI��e�u�EТNSl�_�bi��<�e�(��yT�� �ϭM	v�	t4�� ]�5��ߧ� 4k���nJ���A$��J0�9b���Q���,�� �O�z����	��n�(N�jr�g�NI����O�y/3��E.IjMxEp��KqU����I�!Ow~qAF�O3�R�B��neL	Xޖ�w�-�Pے� �6��b8��N;R���PR$
�������^K9�)�i�S�]�<O,��a���%җ��
�p�}ZK�-(�#N�7l4T��۩�?c O�m-�
�@p4���(Q��[rPq��r����~�ړ}]-e�7?�&�w��펻��
P��ɺ�]��	��^x�Ԉ�t4P��6���&�G��u�o�D�lX�Tա�Ҫ��]W-���FQ�+���O�=|�����[@�f��^�s��PK�	e}�j�4�g�-��d��#��M����[(>s;Pa^PV������GJ�8#e�NS����|���W�]p7���4�ޡg�V�)�>Z���3g��P��P?���>s�s"T�77��۬y�K�T�@z��|����T.7tM�ب�υ��b�M�#ЯƤ���Xϻ��d�M�2����q�J�/v#��k"��F3�q?8L;N��N����o�-O'K�9u�B�) ��H�{,�DS�A�Y_�d?Z�/�"hڀù#�S�oK�o�S���#C;,��h�(�ݨ�|I��Ŋ�������=��U���`.�AG����͓���-�tH$]Z�Ԥ!FV�Jj����dU�"�n	4k3���%V��Lh����JLC�}Zh�K�"|=z���g�Zct�v�C.銈��nE��KS�ǀ����x�7�|� 2=� \	�`e�=1�Y�aSk �E�"���G�gCϞ��TU|i���Fx�G�ʒc��T��1s�����H��a����t��tu˲���Ҫ�2⺝>��ע���.j֛� m���!>\x@|RF��X����ֲ]�jBPע���EÙϗ<������=��oB��냓����G��5Y��[?�_H�5cf7Q�&k`b�n��e���i��I�E�T�$J�7���i���/�~)B�e0��S����-�^=��S��VG����P��`d1Ou�5�e=i~�5xz�1�0����X�JF��^�t��t#p��Q�s�`�V@�&�70Wq��z���~���#e�ѹ	%�C?��na��lFVL�.=��Ԧ��x��Z�w����%A�B�=âܛn�����;"t��~<�	h�x�)ph��%t�$�UD����'8�}�X<�/��v5Y%f�u@"VV"FpV�����|=� �[��v��iIϥ)��"ݓ�+J����|����0E��>�*���mpe��r�G��y�w�Q^�Q�B(R
�3ee*������䮢r|�Jǚ����@��ϻN���j�����v1�Q�e7�n�;�p�cB�r��B�����s�L�")� w&��\&�<�}Z�5}��-5Z
?'u���Jw2�����/6wn��Z���Щg��.XJ�OeփC�q����>�d��?����Z=�ílhw,�ڳL�IJ
��/�[����mG���C =Fn|�Y����j0%��bmtm���P�Y�38ul�_�UL�J&��qYJ@�ꎙ�5���c	G�t�+~�P���)(p5�bH��ϋ1�����Ҽ�.�d��[�l4�K�y����*�=;�����̽�/sc��(�3�IA�2����2��մ��08H��TTc�I��)7'��+GcgZ��Z����Ԫ�3�t�a9�U��!��8�i��,Ｚ�&��%iL�V>J��+TR�x�k�+A�?����"�l*��~s5/|H��� �b�r�c��D�I�b��pi���^Ms1�_ۭ����+�Yx
��F<a�"N��~v�������p�m9ʗy��s�����F�A�_��Y���&H:Q�J�+��挤�6��O����H�=��$����s��OM��$�c���#��~�i���p��}A�9N�bZ���(���2��xxPw^�����ڏ�s���"�~y��~%6u^����l�K~y��n� Ȥ;p��U�E �!�=n6!>Y���F�K4�0~\py5xVJ�z�y�В�&�/�L���Y��ĻH��RV��\�̛]���RqICCr�@-��۰�#���Q:�g�G�����e7�(�����Nd�嘲�;,[�!:#�����0�90�����h��j� �.K�{����T���+2��vyIЬ�����@I4g�~�#� ��>E��G���F%y1�����y�;��f��j@�\]m0�0�t�CI<��O��� ����\s(-K׀O^[�"��ؐ��ꞕ�ö3�4�b�%|��E�8����є�G���s�:[Sz�q���힉�����̩�<�c�̈́�Q1�Z�O��VO�p
�A����>���}��"�C�:� �-�5'<�@'��ͩ���p-��vbt�@���>�G��A7��9�Ra/g�ᶮ�������G�B���;6�ps��	]���&�Vs�S&��Ƭ+]}��^�1�iX�� V#��W��'f�j݅�r�fc�Y7{��d��b�?�b
'�Ld`����"���H�p!�2M��r8�:2f�#��/��TL�>��w�f�9V�<!���{Sfr¶NJ 2��[2��c)�O#����{�����)�k�3v�{�Aw��ȧuߛrF�h}��>!��H�7��X|Ew�/݇�P��)檷p�����\�4�"�.G� �j�Ob}�:c?��mL��/���=���û����!�,l�V�Z�Lb��zK����Ȋ bn���Q��;���Q1��vv�uG����/QZ�x�L�{���P�%t�k9A�!�.�+9?����#3 6�H�J̙�Gu�V�T;�����F�/�`{�7*&���%ǵ�RH�>.4�T�)���P�éO	�Tl7���%݂Y�'���Ӊ=|i)(�z��Lف\�J�9h�k�#1�����3����$��tL��BWRѦg�Z��w�n@�w�X���k��QE�l0�DA27W�c��`��ځAӛ�u��qh��j���=�:�?��|���|I����N�w˗�Y�6��:��d��YtO�?�Q�ON�U�5Wk�I�\U�aN�e.G��4�{��{�F#"|� �^���	��R,ɬy�<#��N~�����ܟ��EWD�3��(�|?	���ܝ��w����0�_Ƞ�x}��c��]�a�� �F	�����:OD-�}t6n7�<���&i��J#��'a#�xO�n}�*�@�뿫��������_�H��ɛ��(��l���� h���E1�lZGXe�_̧8��C��v$KZt�x�����~����&���s'V�X����Dc̮c����q9�V��EY+��(����ʔ�O�L֖p��Ȏ�00��K���u�����q^%��68tO����u�l���I��-�IP	#���Ï�_����iU����8D�ښ@=rk����MYXE����M5�AOλP��AĘ�3eI	<�mf��)��k���䖕.|�"�����"\��أBk�\Yu��>������<xl!1�xUȷ��cp�����Z.���I�g��	*��\�
`y��P��Gz��x{�P[?��z"�P}*%���w?\��<���S��'"��SpP�<��E�=�O�tw���4��]��j�d�3"7�im������H�j4��T����L��I�B�{�	�\�Y��U,����-�QF��p'����/���?E�jQu�p�Rc⽛͏>l�/c0�y��r����2��'n2�v���z(�� g�L�š���T�"6��{��/��h��囻���b�<�a���c�5¶�Y��1�Gb�x߃�m���ls���+�0=���DҢ9M��s�M��*��$ ���8�:��0�2����gW�B�m����˳Y)��驼�?w(�vV�K�ƥ�;�
�����Ӏ�������uBJ	��K����7$����$�aa�!�JԴ8���G �m�`�����ե��S���ʛ��`���\�i��RsR�;��D�q]�b�C:%��ۖy�����(Z�
��!5T@�mm�MI�Q�F����f�0b�=K4���Ini ��V�8�SlR���gB��u�a��]����c�V�B,�	���Cƙ��2�[yW�.-�~�xP��5�(��S�p�.H������'��#ֶ]��bR�A0L�-o�()>�rt��fi��%a�&#���KBi|ُ<�u�j-v�Z,���*U7&�Ⱦe�3w𭦹C �j~��|ش\���t"�L*��<�j(�Tu�L>8fóm��Nj����P;U*�fY�i��_G܃;��Pn���/��ߑ�*�>�IδH��2�4�y�<���
A���p��h�:��:�$\��i����z�yS��z�gRc`z;����|�m�>�i�a�n�1�ǐ��<ȌZ�'I+��#�D�\5�T�~�Zd��eC�#+G�} ��Z]9񀄲	�ɹj����Iן���x�9
@�����h�q�7�"탼MMt�qE���@D��]��7(�fb���Z�㺢v�?o�6�H���X�l'#B�����ݴ��ń3��ҡ���U�!*��&"����)��U�ِ>���*lI�� ���0ayɁT��k��T&���'�����ĸy�r-�lQ�i���6��@���+�&�2 �/�/p�wG�����������؏�>[�j����休�F�?�F`��ɔ,���<C�E	�fq��ձH������1u��N��8s��ȗ�;X���tώJh{�B�l��q�e����;/6j������t�s֝%�����|lH��r$f�/�n�w�T=���b4,�U�tO��$�S���}�����kD��d�� ��dk��;�'�/H��(d]�B�*�r�|�l�n�� Hm�i��˹!��G����Z�b���%(�%�G����Cy�Kã�W�����x^���'��<͔!z���2�dgce����D�'yM ă�����)ة C��A�i^�J��O�`)CO&ފ�P�G���Z�l���6@�E� ~���C
�9�,5f�\�n�����LQbM��%���!Mw���d¾���9>�&G=�u��޽���gĤ|$�C4"��K����M�>�44�ae��x��h��"���;h�����X�D�-^G�u��� �mq�*�4�Xz�ؒ�����\?űZ[���{�XUG/{�}j����c�;����]�J�wn�<��_�<(�<�M#W�oa�N��VI��j����x�\�w������qg�r\�ZQ���\�t�Mύ�F��.*BF�Hh?�Rk�u�����4�����*l�i7Ta�	Z�7��_AL���y�����T����)%�ȡܕ$�񾧿���5HU�
�|h0��o��m��s7*�Riai��>�T=���֔��U:S��xi��Z�	5��yv���X�K��>#�̘z�.��b)r�Z�����o&*o�~�#�.��N���E�ؕ߉�U�oC����Vӊ�������9Z�9�n���5��1U����8�$���'a��z�2�3S�dO���V��<��̜��Ov�-�Jv]ӵ�k����iJ��'B��i�����L$�]4M�	F���������]���t�-F�/Q$e0�ޟ�S�.��3��o��+N�)���`����76v��T����{��A'k:M�$��P�V����E����MA�e{6�scE�eL�IE,�)�b��؎3׏��l��£$�hò+qJ��]���Lv��1��Kx���-�ڬ����3��� �bT������'ki������<���0�#�zL��� s���;6t��L#���ɜ�E�U�]�,y�?�7=�*�h�ak���Cbc�>��g��yz6����Rw��Ve-�dq��a6}u�U�?Hi}����%��m~�IR�=��f��$�Js}�߳Prm��L#H��	4��~(r(���>cA���@����&`�m�E+[�w���!���(f�x�f6Sӷ�,a���FK�,.�æ
�5�8�9cfڲKä$��m1�
YlP)�bQ; ��8�������k���6c�$'vA�&w�0��m��ߏ���O]���3���c� ��I��y�ȵ�����G�;�
���cv.���e'Ƭ�