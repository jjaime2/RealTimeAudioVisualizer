��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E�ﻏ��Aގ�~ބq\�l�1�4QQB��t�
�_�㬃1Iw�$�=�\�:�}Օqգ�$�ZB�h��NS%`2#r�e��c��B��FJ�CH"!��G�D�}�� �5��7��x��n�{��:~{��P���{v�� �I�ZW�컪e�3��hK|�|�k�/�l}��l� 2�3ݳ�����-*Z06Hf�\��eJ�8����鯚�%��d��9��!O�q��(�8H��&���$�ϻ�ʧP�J��:s����f
����U�m���j��75���!��+L����2Za�,|}�燷�N�r;�z�����]����E���"��?��M���2a+ -�踓�~��ҵ��h��N�+���Y�A}W؜Y�0�c��nz�*�Vr���t�
̠a<��!�f`;�������j������Ndx� %R�r�Ap����3��}�)�`u�Ǌ�GO P)��C¡�����[͞�H�,2�$�|��@�ɣ�zS�ҡ�a�=��Y�U��$���� X��5��qX,F��LLS�T�Qde�����o�c�<���ƹ���?���lP�5��!7�U/g����ْ��߮<��g�Q��4��2l��ζ�B���J��Ur��K�c�&c0�j��͂�{u���e�o5t��.8 ��XC5���4�̺�º�bBS�M�^�g�Ō�>�M�f�3�sW���V���L��'������
�XIo���s��8^�H�T����0~��L��2a@�R�!�����d���1��lc(���|$`n�S�BK��,���!_�->-�ԌM�a���*#�v��:�Z�&g�lRl�Y5N�@6v��iLEk��{�,���'���ߐ�P�!:�,E?�c8�3��e�y��tV~N,"�}�<a:J��қf)����Km�F��KFV�E1>ZH�ŝ�kHp�C&��}�dG�L!���R?�{�g׮r�e8q�<j�9�r��U���̱���%�Uɷ�Q�
�d���&�Xv	`�52Ԛ�GZ��������;�|r�`;��J:J,����7��ޜ���%��>�M��+ް鶬12lO2�K�Xl��gQ�`��1�zҸ�4����]��-��v���:����#���.0M���L���:F#1>�{��l%QA*O����ŚJC�=�����s�J��g$cc�ŧ÷_ޘ3�;��)�e�Mk?���ȷ�/�8z9�Z�6PO�c�Ljt��қ��B}o�zX^�'09��I6>-�?NVC��G����;���3�:�(�q�;��]���~Ă4�r5�{U��W䵽W��__N.2蒠�@!��g^x������@w&`����K(��l�5.p��P�Jm�!�py~f5�Q�;�2m���ӿ���Gxφ����T��	��u�F�6����4$Yt���M�C��~<�T�c�������:��� <��fN��k��S��%[g@6a_�5�ׂ�4Zc夹5Όr#쑣�+T�Y����y�%�T��HM�a�֛�<]/ز��:�J����rp��p�/T���=| ��ޙp�}���7sH9�����B�q��,/���<����qP�"�*La�ɝ�m���j����+=v)�����׎6T6�u������&�tf�m@�ޚ?�
�Yv@�}!��Q��֎|h�f5Na�7{{�b�"�p^�<߭ky�%�қGi�BBԹʫz��ȳ����/3f�䜥���ϱ; \��h|e[D$:	ȗk`"��}"b�]�I�h�R����S���I_��S;^mr��g���l�=Il�0��['m4�9�
`�T��\���V���m�����^ޑY��(�.ً���O0�m���Sĥ ���P*������X�߸��
�}�㣽;Sh�X�Ә�){�7;�iw	1
V
1i H���2.ˋ�x���#+�qO�݁�y'�~|/��D���a��>��To�NЌ�f�~��8�����6�u�;RC���L#j�u�g���N k�'yv��C���XL��qFU�~�Rp����.6��������:�Vzxҩ�����YOZb�#�9�C�n\�w��1Qh�0%p�R'=�^����
3��Tqa�Jq'�֫�
h��������H�]�NkH<���L�Z�ˉ�L�(�TX�,�������  ���N��y�?���h�eV�h���J��(XI*�Y*�OG�z�8y�q7�6��޾�ȊK�i��*�voG����`�5$��6UF/�mM�)����[$�6W/�Q�	)�R�Bm��RUS�'�mk���5z�)��^�����nX 8�`*�E�V� `m�������Z���V����5ӝ��sh
�Ɍ�EQw����-��-Y�y��s�1E&#��lbD�X1cKej�i4��-�&����ٵ����+^���ti��s�uf4�J�8�����+��%���fF���I�e�Q'���wue7�˱G1��p�&��Y�T��v��@��K ��2� �r�V�_�8��㲙U�O�K��!�i��;���y�Х�4ϋ���,m��ڠJ�@Yv���ʴ��;�=a����"(�#0 p�6^}-j��Xb�}�~q��.�x,N��kS��cX�t{ۆ9�����kBϊ��y�-�ʻ�	��SzQj��u�FL������A؋VTwsnx0�5s�)��0���J��d�w&k5��R���";�D�)�G!cid^s��l]�D�+ʂ���g]�?���y4�HT�P�v3���s@/o����y6K.CDX�x�����_J�(��8]r���ӯ0��/r�^�}`).�.����x�8,�y,��Łi4w�6�u�ҧ����	"5���\,���]X.F:��;��`;SUM���n��Z<��t����YXܨ����{�^%��$l�X���J	N�Hf)��,yI5j��X��Myf���"��ۑ�`^�@R¥�-����&B��+̱i0f�#��D��>��8!?��Z�S^9�&�>��"�b����L��.�+�o����>�5)j���Wim_������Vks�ط �6m����"�y�9g��V�D��>C��h3T���r�rN��ʜ�-�ښ�/SLƪɠ̣Ѧ���|_�M3q�e�)o.�ó,���.�5����S��&�pZX���w�)�̀8�[<J���n`��\"�����fd�dQ@ ��!���������d8�����$c	�$d�Ϋ�����e�wn�5��d�>�i�8�A��5��As%J�KTY�?�aU�X����1��a�����QAR���܁r�V��X���`��eÚ��77MM�6�� ȇ=���O �G�s$�e���h� pk����y���;�1�c�C:�<��Ǳ�h=iu�!��[�a|�Y��r����k uR .�B��To��dC��N©t����s!� L�� $�,o����m�\U]�Ө�h[�)�\,�9�ȶ���#�ܞ�8���%�`9L�\5r������+�]�X��a\�V��sɤ��q�N4��>6��i[!��>ɋVR�Ӛ�n�3}�g"���%��Dc��wF�����Z��SyX�a�)C��=x{�P3.��=�f�.E���w��D���q���Ԕr[fj0����P���x���	J�6
�lV�Ě�h\ ��h�f:���64���R�J��jHۤw��M��e�]ӓ �C��b�W�0��mZKi�s���|3E�|>�[����>ua��%��h	:-,�u���\mw�}^��:+fm�;6#v�b!����	���r|Q��ީ}Ƈ��%������Mu��aέf���i����=q�ѩ��_�rC��/�����>�@�ם|c�x~;��������H9����)������O�����b�<􎁋F��ޫ^��+5�f�-�>�b.�iIb|t�=��&��&��y�Kf��$C1S���C�G��73T��{�dr���D�e��?�X 5�{�h��v:�� ��PyF_�7��ǁNx���/�<�3NZ�򎭥d±��|��V��s��A`�X/�xL��M����ň�9�hD�<�j�������E�ڿ�� �4����Y��r�'�s�|��A����N���B�,Ll���-�h�,sa��à�p<4��Ja�öYk޴L���Ä��m�j��%� ?�851�qJW�O6�w$��C_�Ƿ]_��`p��YSN��Cv���y��*�hdr�֡յ9���SR.�@N�/�9�����ߨ.�7w�l�QCW���`|�D_�:��䐵����"@�Z�T�n�T+���"�s��	aj߬� ;O���3���w.K6OXê%		����Xiԩ�մ��G����@��,I�O�8|�4�iԆ���/Vv��ᘇ~}���x�A�c�"���pq��}���&h���k��o�iQﺫ���8�r���&s>�fwWT�u���&o���0~����X��� ��������vae��F3�w�*WNۡ@	R�&��eB�h[?G�0��� b�^�+1�7#��h�v"��-@}%���֦_��M�lI�>��X�gЂ����)*	�Z��\�s�6Չl���-5�������ܭ�v�1E�ꯗ��f � �e��ӣƪ{6[�I�j�F^G/�V��%7Wq+�ҹLH4��f�bbS�PQ0?��q}�_��dF��T�A���^��m�.��Y�dį��@�HGY�M�zD��Z�Us�� �ab%�"��Fn����E�h��,S3Pk���i5hL�4��}g0���>�#"g6�k �E?fV>౬�q���ī��/+˪h����L@���t\q+̤Z�?�3|�&,9!��_����y�u�|ų������όS�L4YJ�N�_3�7����ْu���Ō����V}�0�b$_���C�E�nHԶx���>O�,���L�Ư5Đ�+�6P@��ÎfϒTJ���x~bN�1�Ĉ�?��Ӓ�>d�v�2k�-���Qݯ���.N�hb�����:�)��Se/��f�c:�ui�+H�Xu������&�W:`�Le��۽-���?m;�6D�1tG�%��_�(��G�%�?��A��������y #X��9���R"6$~ !�I:����V3����xX��hHC�ǮY�
��}K����XEf�֦��  ���h{���Pdu}	�d���z$�Q���7��9���TY )RW�1�衔����gm����u��FƦ��-�n��͒�	��b0/YD[Ǵ�^��]FX��s�U>�ٵ�pk�������L���}���i���^."g���^�T��F�˘A��\x�k?��O�e.m�+λH�]"�Q��'Y>�u��\��5u9�$����j��
-�K���}m�O�ڜ�-I6'�?�������
�I$WD�Qdhq����&�UI`Q�@��T��������!ڒ��r��l(4�$�h{&q��k�C��C4w����k[[�Psg��������{�����##��ޔz,;u�e}�:�{`8s�$K!���"ဗ΁���W����r���Z'��K�<�V~~W��Spi�{E�2W�J�0�ERp�{jR�2:��u��?��H��\�0UuC�+H��4�����,c��g�K1+G�)D�)a��2�eo*��|�yjd
��b�`ZBAސj�$����l����:}1�4�/h2s��F\q�}����[� �&|"]y�0�X���3�T�;�k��1�ú���Ή����!�.Ū#�t�<�B@h?wι�+r�d�@ז}
n��;�Vn�v�ǲ(ZK�pB��J�P����D泙��UC��iI.]!q��=㵃Ir�5��]�'j�Ki3�=���d6hx`�Y�ѿw�]f�!����r?�