��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#��R�C(>�-|+����J;���5ǔ8#.5Ⱥ�`0���Ny,�iOK�պih�W���?$���!��p�n�d�v�O ��E��C��V͐+@�v#z��O-ћ)��[����:�-�+��K�K�ڍ�=[�!S���7��"5��h/��S���v���$^8&A������Y͹D��&�σ�ʠi|�AN�x"zO��fRTy�������y�M��e	���xyw�l���@�H5@���c'�-g���pDO��d1��0�Cl�r��q��� GdO��Nz+�t"b�iI���Q��1����t0�/�#�`'w�,���?��'f:n��Ǉ�F�o]����}����_?k ���L'���싔�F(6�-���C�R�{�U9�:��XeP��j���T��.=�GC2w�͑���Q_j��d쯕]Ӊl�he�I��cS%���S��8)yM��pW��W��?�3K)3����2��4�~)��˾s|���{GdXm�z|��k�����U��E���b6�o��epY��	�$R�.�
F9>�/�r|��w�n��X���xci!�	�i�&s6,1s���IN����b�����n��`C,����F�o�vd��<q�l�¥�����*�e&`�uo��S%O�p|>WE5�P��_��p"��^I�|N2`�锭��]��VB�����>�W���G MD�&�c��L��k����g�jĩ3��f��&��y<�ڦ�W��I���fg_*�F���^����_#)Sƅ�J>N�?#.6��:e����G�=!���z�X�C�q�EXG)�.JR�=�B�
AS��豌���,����@o+lwQ���,��ONnoiv�����#��i�/(y/U���^B�Z�7��
�6U�mX	��F��ku��p3`����;Ip�%8�[�Vk4�j��,B����D4��������[�`�����jF�
���y��ƀ���e v㼱���ٷ�ا�r�l��W�0l�,���$�ti�P�<����s3�4^��9zx����}�����:��i5yؑ�� ���������1q�W�����fI ��ώw���c�E���%nrq�Pd]���c̨4�3)�,�<���-Q5��*�.��r	c��;n��*����Z5��`-���U��;���;��}�tp6q]?+'�s4;��/-�<�PŃL��I���&�+V%���0\�I�h�����9+�;��/@�;z��Й��k�s��򵘝t1���������i��v��cL���5�� ���w��Rʺ��x;Rq
��_���H���
�@�����o8 ���!���m�[�뺴�;��}��!�ZGs��o�[�~%dt�����N�WX�kq��Ն�j���j M <���}�a��}{���n��Sn�q�o���+��`HH1�t(^�`�@\�u�����%w��H^<Y������]K��.���ݝx�DY��7���j�:¢�J�D^��0JGH�*�]�=U�i���,�f p�c]I�ɼ��9�dI�,�m֤�W��yɱ�m�!�qJbp|��nD2F:�o ;�����8�Xt���K��!�* �i�f������[+���b�&�� �ځ���U���b+���t�m#�����,�Y~��t��#���R�`��"��x�;�����A|�d"�� �!I��jP�m?��</J���h�\|�6�6��.�� 1����h�\�f�\���fO`2�T���%�/�0� ���m��KI��2�F�(��CН3���[��#�}���s�Q�:�f�^�Zb�OԳ-��,��:KD�v}7�-&0�8���HH����knՠ���_�7�,V�8';�Z���
��IwH�*NsZ(s�h(�)V���MC�+� �����]`<��:�K�n/s����e��ՙ�wZ�8)��Gh���u�h���}�U��Q1��y T���V�
������{�;F_��Ԫ�r���4y��j7[�9xq�Dv}P^K�
��i^u|uo��X���1�F�sĻ|@6���Y���5h(^ܼ|���.>H�"	��\^��{�|�B�H�G&�A���W0�OzJX�|�}���� �7.`|64V���kC2]aB�>�e\xL݊�!K�����N����Ⰵ�Mo0��>�Ř�~ۊ��\����J ��!L��C3`"�2^.Q H�>F\�NaOYɴ�dԁ���5ʶ$��qX)`b�{� �:�$�I"�=q�J#��|ոNsb�y�H��߳:!Og�)�4�^�)�jRv�jA	�g䛢}��Cx� �E��P1V�(?��� ��X�ux��}��%�io��f�7s��u�aJ�)B?4>QV�����^~�Q�s���d��)i{:��"�������V*�Q9j6_�6����é-K{���ʳ{hE;L�y�ӆH솎E��?j�8���G���m�l~[۞$����_=vfMyjze�W�w2��K��g���o�Y.�b2+�.�F�q��}��\�m�
�����J�0z6�Cz\�����v���Ʒ\����ص^�,M\��>� �1N�+�}��4}��Z�?N?��Z�xT����L�P�0����d=�W9L�bW���f���zо�]���I��� �-k�N��`�沑���1�����	U�����p�rV&�Կ��MŰ���U��& )��r�aQ����\��*�Ǘ��o� w�qu�D��� 8�L�6���I����+`�<��~ u�u��x=W�+���qzۥ���1pb����O��"�A[`�x�w��e����=QıB��+���$��dK�c)� ��8u��+~6�(\~r"dV�E�{�����ɒ��>vB$�Ww��<j
3�y4 nT�Ve��?��m����g��	р��";����{)P$W��Oʬ��i��^�Aw�7#�����{���)+���ڲ_��1���ڲ����d/g��
Ā�\�U��������Q�<��{{!c˓()���v����;�y4�ͼ��Y��Dl�[Z����g�ε�$=��,B�����0�[�"@�+�j���m, +��dD;�{��U�m6q2�����n�r%���R A�v�����D<k�XD��#�bOq\��ε|�I�L�iə�! �Glk�+�>�c�l�۱��H.�i�x���T�]и�O�*h���6�?�е̳�M$3�W��:�<�Q2W��7������u<! �"=u�W�3pV fށ�*�XeЃA��hr�$)��=���t�ɻӊ�ESl���\5"��i&�+�f9���2��ɒ�&ފ�{]���e��l˶�~Ijx�Q��F�';ސ�i��0�]���:*�� 7q�7�q�s#&jKP)ϴ����v����&qa����R(��tX���h��4ã��&p{��z�(���;�+VF��"X���r��#���E��SӸ ��u_��	�`5#'��	�;ƹ�����q'#�η/���ڥ��e�&�2a�tݮs����:ų70��0�n�$�"���;��տ��W�H�O\���>�,f�]Ẳ!Z��{3_�n�\�q}.�B��8й�j�	z4�C��Ї�a�BH.�̯�W�iQ��D����L}�](�TD�?k���IĒ��hjz�����-ɢO �U�N�٨16\��E��Y}�{b�D���	���7rB9����G��JY���)�a���~Z�4��H��8D�A�Wl)T��[5ͣ �4����3�jp��������]�Ͻj��,��O0��bd<�䨌�ٮu:�1���q���V��2�b ��e
����2���ph�+��ܥB�aH�5�F��sO�