��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D ��(w����E��}�U.��K0��m�A�x�����m]�ǟ�������"m81T�A�q��z���7��M����~�`�]����9�Q��qۘ�C��
�'�//T!�ѾbA���sq�]��[����A9���:��+�<��s�A<����?����C��A�5��i�NV�V}�������X�R�R�=���\H�2ŝ�`tw��	��v4(BT�����:F�Sݼ%�+�=�1a�M���ދZ��q�7�/K���:	��&�_�V�V!.6?(S��o=��m�4��X3ϥ	�6��ĸ�����&����2h�� �la�|U������F����gf:a2�SFP;�� �8 E�:��z�6&��A��K|��]�1c��NX���UBO%l(	`Lڱ�/�sӏ?�JG0�BV}����p�S�QF0��B��P�0��a�h�yx������C��@���L��Q�*;+ƫUz�	��.za�����9u�8��}_a��-�����/�&�Jl��ϳ0��V�n�	�J���j5c�����<����Z�6)\��+��`��%t"�6웺��)d�]c)���m���k�������S���ڬ��j�~?��A������d�� T�\�K���k�0�7�߫<��g�\h�J<n�@!BK/o�*�[�G����k�<\��T��ْ���b�O�h\������s��cgo��ю$� .�:un�j穀;{uܣhС�Ov�(z�3eW��=�>�k�1��
��Aw+�r�I�&��aLG �x�p)�n�����f�}�h4�G�]҄iĦQ�@��ٴ	��XpR1Ƿ.�ƅ����1�i�eď���V@k���gئ2��m���זcR�B��1��ޡ2�{/����d�~�Pd:�l�������o��^6QJ�4�������H�����r�a�j��Q�o��F{�}��t�GI?��A�n�X(r�/����D�/ɷg���L��o�j�(�<��G!��2+㒠��)����̿Vq��q�U@/��-�����(�� Q�v�# ����� O�o��Q��2>K4�{�r���8;��I��&%T_Ă�5|�%\�r I��P��nO��d�� �KS^�������do���
�P��F�ձ]��T@�������ih�[��-�k��]F�ߙٌ�
©͚�f!�=%���d�D�u��ۜ���CS[�����9:̢�yQ` �Q�w	�67��p�cVۆ�},�)q��Ƒ�k��dE佺�p�[�@Ձc�\h"��#`�ܜl\�!TN��R V�_�!��{�D�,j�uP6�q�IH]�>��Αw8@̌\^5u�j�$�Cv^�W�7���@��Ǭ`�E�R��M�؟�������0�qb3\]��uJ��*��)l*ױt�J>8�
�>�3,�D<��l�&�m�0^�6b�ΧC�;�&����45�E��/�/��^4���_��W�=ی�~&Tϒ��<�5�7�"�<[O���6�^��hQ}<p9�_,]*�x[�"?u�.0��[f_38˭�ߪ�O ��C�z�#�`��ޒ|�����7N�1���$�����;Wb���
�RuN�ay��x�0&�l$�q[/�'�D
+��Ecл�o��դ"EE_��'��=j�$���'�`4EH����yuWs���`������e�!MF�A7��7�):��n������o�c<2�Ci�-��y���װN�Z���wd��i>�!@�YX&�z�tJʴ��ѐ���Q�~<'h������+t��Dܛ�L��f��܃���A�R����A�8�`��A�h3��ڡ�m"Q�ļ얺�u�|�)r��%ћ��{��h��\��9[������K�����G=��]���H�ev����OW��SH��ꈀ���'�ؕ��]�ߑ$��I�^�h���㱆;ǡ �KՃ_S�a92["�zKJ!��{A9�B�^D���U�^h8*��'[�����S��m�Vv6�rD0QJ�TJ��Pۈ�j�Z���agh��@�F$oE9
�{��FPKRY�x0���h�?�b��l4�5��c�N�CR�I�4н]udʌ�Mt�
Ԭe"L  Y���]��D��9��&; �<}˱�(͌+�suE���(\�.y*bgR:�&������{!�\+�֖���>{�7m�mrg��wD3)������C�PpoJ�|Z���K�]Kkw�� ���_���m��w�!?g�ŭ"H4*⬆��W}���f�]�0�
N�۰��h���k$M�-1�f� ��BO��=&0�����di����Xl-����d����T"c�_{:��:�Ĳ��r����Yu�WpIpS�LEM�
R7��_�״衎�/>w��,���?��R	�3f��Po"M��'������>��s#�?,�t�|��q{��Z�ҙ"Xw�%aZGçS/���܏���2�S"D�@'�D��)�x)yl��W-omv7��\ZpӲ}� �T��*2W:��/�3J��f�*��M��C����w��0�A�M��Ho�u����x���d*O��8���h�p���?�`�Wᴫ���S<�>T�b�������E�w}0��ǿRbP�>1&�n���Nf�|>be��`EO}�)5��CV?�Z���>[��Z�c�E�?r�څN��\N�؟�� t��+�?=H_�����ݽ
 !�n��k�"#������Q2ƌV���i���}��æ��mo��|�M�?J$�[��3��[A��+�'�e̹���2��#G1��G����g�`���?JG<Ӑ��Y[�ST��¡K��t9�Z ����34a]�xy@��M�:�$|�qڋ	� )N�2q�52�89(:L�.M�*��*��ٿ�ˬ���lNL�j�6�{+FC!��֙�;c,�%eu^~��DR��(h�������ܒ�i��%%��=/U�x�ƹ��7�{�o�QQ�d9W�D����
�����w�X��0�`B�n�5�V���E(1�������RBVcv�������Ӹ��A�)�M�[]�9������������s��d�[h���SW�x�,^���&�k�ɍ�:\�bvzH�6,	wj7�n��fdۛ�����������@���%d7��P�ޡ|�����4��2M��h�򯕶
qc�[���ym��x"n	�(p��K�ڕ|�_�@m~���p)�bj61"�2i�B=z����Iؓ��W��q�mV��|���ҷ�덠jW52Q3iЄd�����<��A��u�����1
S�1���t�Z�h��~�ϖ�e����_x������� ��+_*�0_����V�G�2G�	��w�
��vλ���Q�Wp�c���Q�x�>��"�_5(-/���:F��N��;��9���5�F�[k�Vjt`����3�I0����x��޾��������� �SD�nz�^�ŘSv��Ɖ	%��8�����F\�W�b�K�m�j/������'&1�?ۻK�ef�QSE�jeC�n���$e�8I�R�9��J=s�(@z�����b��gפ��J���JQ����F#]K�6齚V?�����+zB�oY�^��{�S�Cx��3���+��x"O�����Ⱥ��yHo1�̴�KƹV7U�����������k�/[��6�м���elx��5��&`!@h�f�<���}hʀv�UQ���)�
jM_��i߅�bՄxG�
^�(��<Z�<��&�r��r�]���=)GT�qϬÚy��4�U�?�oH��
dXp�]7^"	>�����)���r��S��r�34�L�9h�]y�����2�R��JT�cݨXq�&͈ �Ӏ$�������KnVq��1�aV1K|FQ�fY�9���q���O�6��t�O�R��'���tħ�Э���xQ J!�����0�bu��Ӭ��<�ʖ�{B�VX�G����~�]�qM������z ��m3}^fLL!b�s#�N����
g�*j��(�:k��0�&�;8?��>��~�:L~��S���P�ӈHL�ni�[�MCX�|�����Z,V��R�#������Ng&q�?�9։�6� ώ��2���v�R�P�郎��UX�Ep]�q9H�P=a�I(>	����ZQ6.�� f����o�$`�E����%K�!����Y9��b1�q\�`|��V\�b�E�~^,қ%�BМ�7�'���Oc��O0JϪ2�0io���� �����J�((��:�ϵ=;)��i�'��I��/X�b/U��1DM��Xm���淟Wv�^��J�X��@��),ڥ��o���7�u���)�������2i`�Η����I��M��@��e:{��#��{"�q+1��4d�C�I�+&Z=P|��i�Tf:ܾ̓�����bK٩�"˶N?�-�X1�_2���v��\�
���G��xax�ӓ�s���Ԧ��g�A���T(r�8mLmʯ�Eժ�-Dń�\�\�<h,R-����[G�W�[��3L^{�<�D�>j���j<=��u�QD�������&PC�,��V�W5�K'��M�
��*lpAI��Z��e���m�I�w�ٜ��w�]���'�y3�x���8F.��}�T�é��W�xZ�������}�����R���:�C�ҹ�L8�6>E��7c� .��X��*�����>%y�4�8嫶�^~F��d��*�ϓ8�<��J���.�D���s����ɞ�OґXH�T�f$��P5*{@���^��'��n�U�ʖґV[��F��:�/�Ϙ	A��9�y�˭@wtS֫�~\ė����V+n6���)�������¾	L�vL�i �>'m}� ���]��T�����(M�_.E��3�$L�)	�n�_PI�~B�0CQuT�?�*�b�뿓�e�7�n�!�<J!(�DuS�̵��> �N_�;�CȴsRQ,�3�D>i>�SٶUN˂*�'�k��v�Bh�ș#�p���t����RK b�7-���(%���X����MA�<,Ӥ�A�R��)�#></yIV�OE�ɻ��(\�K��1lH����4i���nH��nx��� T:+3�s�G�ċ0���K�S��	�>d���\�"�i�*)��G_➪�	U���"ah��A��"��Bh��_���C�^�2�G�JP�����]��y�M{��Ɔ<���.�_�|P�O�����j��]fzIa/�v<�q�[[e�Aq�AEM8^��(��M�	CO�T�<��FMK�����*�Q�![���O�%�J��)9{�Z>j(f�Zd�����+=��<!�eI�TY[��2�6Is(����燴^�ꋗ�AzRn\��
�"�s��4jݩ�/�fQl o&=D�18���HJ�W�A�H�ޘ^/T�sO��Q}ԭ��Jjv��9�>�|,>�dOs"�\�	��d�A�8Bcla�eW	�ªrb�� ��A�7����e���.���v��������Vz�X2�5s���P���D�ra"���W�u�;3�.[�$�jt��F��.P��yу����W�����p�`a�(Fw�-�zl��aTb6�էQ@�E]�J��)la���ݝ�}nqX�����!��:�{�`ĕ¡�,�I�� �ž���VU͞���;#G�Z
�>5��$#z��>U����z�`y��p�]:�@!r�&�>c�4���I6��9)���D�f8�uÇ����F�J=`�5-e��d:�0͇.�#gVn����5�Xܓ��*�1�_>:H����,��&�m^�����Ls�g��O����Ν��k�̐�h�e���,;R�$RWPWQb�xQ�ӧ���U�c���i]*�D��,1B0�j����jb?M���-���pؼ�MZ�5�P��O�ֳلq%<$�����1>�^]��+Z�]�qn���Q�h�m�m4�[ꖏ}I�SC|M�k�l:y9�q֙���h�O��n�o�i����|e J]m�(���g��)ogV!ӄ�W�0�{0o,�rQ]�R&ǰ�����TFQh�b�;�||�����
Ф'n��$Z�Q���$>vV$_��g&z�'}m���4�G���7�V,MP�Q��(���s>gB6����߫�=;�
�8T��/_�َ���v����QW[� �g�;~�5G��|�(�5"jT9d�5�u3\xWx؝��R|�P������1w�)vE�Fr�xPv{��7$jq���ȷ�V��L��
����)�A��&�Sq�
�wXG� Z�a�+��X��A�L����D���H��iŦK�޷AҤ�0�
yyD�>g0۵��Dh�^�]A�j���6=�%4k�)Z��Ο~������׹
�r
BJA^����%�!��ғ3�����M�hF��|͕�g�{�F����in�1���i�O�Y|�����	����Cd���׻��~d�¹Ƈ�i�8H�ri\��A���s�4;��I~BKN�`��|�h�a5mҼ�����y�ʷ�<ō��7k��"TB|5�ѳ���/��VH�A��oM(�*/<�~L�#�)����0I�r��G1�A���,h�AhKʂ�N��&���D��3��V����2	y�Ącs�{@��Ԡ�Ӈ���O������Oʇ�f"�M�rM��%U��Jh�xSN��:��ۣ���W�M�$��[p�?+��='��45B��}G�0�Invs�"�����w}� gD4�i�iז++LՓ)����3���G^�o(��V=��G��E�G�]��*Ɋ"~���?�^����bU�\�E5#E�8h�d�0l|�E��)����q���O29��f��jl���v��w��>�.�K�1���-� �@�������7K��ꌫx}��f�z�k KE[��J�}��
jV��
?��vA'ms���p|ʥ������)@�c�= �6���i�d���AU�E��p�9f�&ʚ���k�Q�+Ü�:tlL;����_D+ ����L����X�1�\�����M]$*%�0���u�%8^�,	�Sż@,!Y��ԍ�4�J�\�����fzL�I��R��qN��&P}N͞Wm�ҮOJm�����m-�Z#�M�,��	_Q0`	�L��1A|[��G3���:hX�Ҍ|N�Ff&لO�w�ax���w����4W5�S�$lnG��6�!� ��\��̍���h�QiP�۫��'O`��8�Fz�ү��x:Z�8��dԱ%���&;B�,��ϒXa�*]I�PNP�������������s�/�Emfܮ�AI�IN;^����d�����a?��@A��Z9U��55����(\��p�fz�HJ����O�FJ��Ȣ`�<�D��`r����d���R� �K���BC�h��J�b��x�+k�N2�ze6�؀�}j�!~��Q�.�(@�i�F�{�7�
O��*L���)UF��s��R�+����{�)K����ъa���U�=�lE>��hZu�뭸ڦ��>�7:f�@E.<'��f�2 W
j�GH#����tK��j7�B`|����!��H0J��l��\�t�נ�v�I�K��>�u<=�⻭��[�";��%��2�R�����Q�2�~�rC�A
Q�ip����-C�m���z�V*�`H��i=� ���:'u��:?���.��N�f�,BZj1�8��G$ 3�)���2����W��7��/aМ�n��Va�7:C+X��~�9Ѳ��� M�k.��3gE�w!���Pt���
d�CS�yE]�:ۯ����v�q �ײ*��H���7���E�ȥon �L }Ƌ�M�ף�ӵ6]�0r$���n;8(�۾<h�������1��62..^,��^`7A�S�����ƌ%fh롚8�"  X�m#4�X�|�u�< �0 �Tƶ�IZ<��h�u+�l�22):?�C.�b�u�� �1���o>
ET���t������k6V��uf�s	:��e�����|�����#�"x��şo�@���ҧ��A~�ԩ�!�]=Ǯ˙��ɠ�:��,���1�+V�/�w�X`h�.���XAXM��s�GҞruu�24C�*2g�5����3~���*�����������yL\���d5�TA��1i�	�����_�z6%٥7����C��aɐ�1��W�bʫ�%�t�c��X��=�&��M���/#&tÏ�p�78�4R��Y@�N�&���[vG��G��SA@�a� �j�&��= �9�4�p�: ����Z���"e�� ����qe�J@ �v�q)i<m&&�73���T�c�w��u��[��ƅbx������kn��4�9z�ѭu!�w��޵q���k?g6jW�\�r8I&����O���vu�'@6�?�D.�{��b/�_�����:$�xT���GS���Y-)�j=�J��2W(�
��Q��饅>�����[����dq��JF��Io�?����M�(o/fY�sԺ>U�1��|�|w�H/L�&R�c:>�/�������7�[�u���$O����*m�`�/�	%�:`��i���+rӕ~T	���_~eS�jhwn������s�k_� 3'~��Â5�ZMo)0���y	���aen�?0?�;���di�5iE����(X�[�mа�j9����W�W��l��8e�&%1*t�(��w�B]C 2�z![�B�Y�i���]A��^?g�="�M8r䢎"@�7+��鼻�i�U�ۈyj`��8�i�_ ʉ���'Y�I�)�+�b�*Gh생��n������������ �|	Ql��Ŵ�ZC����wqf&P=�X��-�2����`l�p��A�cm��8��e��$	a��|@͟ъ���6���X��db:�c��ܗ�['@�'Ө8�YYH�&�w,�C���D�N_)��ܢ �n�m˛�l��h�*�-��[����?R����-�=X�-+WH�����r�~�L���spO H���H
� �p�GF=�0?R�Xs�J�[���r�k�$ô[i^�(q��b6�<լ�S#�5]L�ɫG��I�p�8��+ԧ�些����Yđ��4@N�F��j��:���?�T��	�+tA
]�X�{Ĺr���_���kwO]�U~���Ǻ�n+�,M���N`k��4h)��ҍ���ך�7BD�E�@<�^�˸b������4�����@�'���=�cF����O��4ݗ��"k������9��s<:Hal�L��%�h6�%�G�0q�T���U�?�\*rb(Ĩ;>M�_�5s|?����Kc���t�m7ص��#�_Y�$w����y�hU	�*4r�]z���1��O+B7���ξY5[�m����v�O�(B�	�hmHJ���6f�n��:^���2pv�O�moa���G?bN��"9�~�� ���E��b�L�wv��R���ʄt�[�,�\Վ��Sͷ�eJ�5rj" X�{���r2h3����:X@M�M�Ө
��O�a+�n(7�Z �I!�iOr~�eo��O��_��ᰛ����C���c�F@�Ұ���2��S|K��o�@���xNK�ٵ�e�l%ZZc	��i��������y�"�h�=JMX�"+IsD�t�ob*p���y�W���H���V�>�]�o��Cc�2_����"���kyfW�l�tct0�'���%��r��KK@$@���3Nb����B�@�9��񚝨���Cx�A�+��U}DA�%M� +/
w��{&��o}�t���3���i�&������^�|���Щ-���q|8�޴�GLR�������0��_��s��?��3f�wQ�ֵ����wN��4o�p�!��)�P�m�9�J�貦�Sz��"ǲ�X�)��7��&6��b��8ܫT%7LV5�!�n~�W�e���mi^�ȶ�Fm�^�^˿V%�HkЭ+�7G:<"��ѻJᗉ����E��bi�\���g���Q2i�	�CK7d�_6%*��񆊾q[� �˛s��3U
����}Ë��0,259��gh�H�'�c�|��6`[̛�����c�vb.�t�ק���f��Wʉ���m��O���F�\��h636-}09���j$�:3�XŞ��%�{j� M�ulԯ(�]�3w�^��lMYid�eNt�v���GU�5��\>|`-���pJh�S!��d���D�Z���M��3ycD�Py0�]7k��Y��:[�w�K�5z�"��9�\��U\�G�Y,쇢
!�k\��݂;\5�0���]Y�4ކgEխ��z�	���T��C~���98A��1�|����zbs-��7�MF�P�a=`�݈����`:�L���� 2��>���pяDsN�.5ڦgL�.�J@J���c�+͊ŗu��I=��瓱�_��൚"ڕ`�bÎO����&zE����p��)��6>E�	��_���2����nzAWY�5�Q�O�4k��[k�$���-+`�4�&Ƌ������6a��t��.�@S�ma݅��k�c��ϧ>[�G��ZE�+`ſ��.Q���oglYˎ��b�oޢ�f����<���0����g]��^of,�2���F	w�%��o٧����H �=�NʦԫDB�x��K���I���^�6е�;��Pz@��m��V-�V�V"����q�O��nä�f~�˗UuфSd�����z�)�S����,-ς(�-��(�m�`�[�g��ON�M`,O��j���N
��d`خ�Ͻ��/� �����`=e�v}�]��9����C�i����gؿ<��4���σ��R�ǵ�+_�I�$Y��#rsǁ_���޿�J��u�/�P'7�A��M�曌V8@>�ވ]x�Иo��t��2�1-���5pW��gʹ��9���!Կ�
�4hb�6LXB$�؋"�t����.c�u����u�n�}wGy�gヮG��z]2L��I�{b�Q��S�d��o{G�?e_
pU�Oe�h\m��Y@�J����=�=��ӕ���D����PFw�Ɵ�9[�k��F���_�����l*<��U������N�P��	���)���z�)q-�����h,�y:�ҫQ�8R�� ���%�Ӯ�Y���k�O�TC��kV���[JW��m��|MxFJ�3R�#��';#B�ߪ,7Ғ��q3�<�E��*x�î�����?�K�������v-vJ~W�T`��DC)� �+����r���//�bM�ͳ���`}�0����#�hQ㈻wm���V}����}x�9jI��s6d�g��9��8^bԬ��:��M�q�7���5��80V�q�d��='���A�k�k�Ӫ(�� bRɪ��l�s��]��ך�u������H��&��VT��N��������3�x�X#9�e���a�Ϥ��z53�m�U[���1����>ljG�48�F"�/�2
~�2�T�F�d ]G1�G}��IiWZ�l��B�|�����$��\�J�E�Cj��䣯��c��oĐ��ۤ^���1������g�Jqw\
wį�Bo���(C���S�s�Ƞ�y��b1�64�W{щ8��xc�a�1��"Jȍȸ��t������'���E9p\�����>A�b�꺜@���ٱ�AH̺������Yd�r_�u;챱���Pt�Pz{����*�ӷ?t���=	���,r��y>�Nw�a�8p�Y���
��A1��Jy�(=S���`J��);�ƗS��T'�9ݛӽ;�v��D��\��)ˋ��y�v�2,���m�,���W!~8��|�~�١�������x�u���WĻ�۠/��qA|ӭ����A����5t��%�S��H���+���U���ˮ��F�7��=s��σk���O�����D��wVR=��xq*�wv�2��fo9]�����򘩥2R���Qj]�j�*����D#ό��\lf(��U.��  v².�,��%�-���V��j��{BO;�L�d���_�Sə(�M@��rn�i��
^���a�����a�bs���4�{@���0��<6w�����{�,_]f5k���;����M�Gk{_�&dTJ�<i�
�����E��$��ޭ�D[�"�p���=u7ǐPF�@�)�]*�]˫�����_=YH�^���d�-�i��]�#bP��o�s�`�	�T�~}ܗz�u��J �����"�n��e���|x�2�7�q��ch�\�h�j5ɷw6��)�|��H�SS|a���
���m���wB#�(��a�;���#u�a�5�����w.@�G� Y��j���ᛯ�,�
`&�=��13}�?�V�I�=�M�˭�5"���#��I�r���T,[�n�~ޤ�c���w�9=��ż�\E���R�T@I�2��
�tvO?8�<�dqyN���<��Laf�ct�3���fgm��3�o���2O���}w��Az��c�����Jk�t���;l� �h<j��� ������js-]��wo�������5��w���1�"W��B2�~m�g��C{��s D��8���P-!U��&��i�sk��ߕu��o��3����sM�~] �H c��ū��Ѻʿ���=�-��� ~%�fE�g�UdQ�"#�O���n���[��*�&�= ��ўB� \��.����a�p���t��(��wxAiv�TD-20���pP�,�I���+@��M����J� Xo� b�Rm�5A��0;����0��CP۸>-�,R�9�)��ND�
���~"в��J��Of�'x�V���B�"�|!m���B��k�DZ�_�#�c�ڱ?=_�^O+��#���⏾$���ն��&陰7�����Mc���[J����~����d>f@]F�	sey���'��6MMB�3�v=n����s?�w����2�����R.���<f�~<�Q�Z���մ�bp��%E����9��v�8h�(��}q2��G�_W(�[H��e#8Ԭv��L�H�MC�P�`1YyF�r�C�zSB�������X�E�J�O�z�͵<���J���@N����a̛���Y�(��*����U��Y��̝��"2ض�<K3�?AP/%��$��w7��������rn��ַ�˼o�͟�1�Z�KG�<���'b�x�<��ѿ����?}��}�V���;��b�tX�7+�\p�����o�n �Q
��\���7H���Y�U�����~3��Y)���N�u�8�op�OU����#䞡���,X�9����~�G�m���ufw�k�P� ߵ�61�u�zS)w��aN(0!�ei�Cq!���E %�1p9/��S���l�:��`�&ت����v*GФQn�J�$�K��<�����ga�|.�N��Q��=�p��ot/���b2y����� ����)��U��rV���#7��93�J�1L���+l5���l� `�+�(f�i�Mh�$ʑ�D*�J�?A���Ŭ�guV�fŭ�Ԟ���s%65��/I�`�;=dW���LM�tN��J"H/;�>õ	G�:y��!P�`���7��_9E|.KE �@$o�Fv
USh��9	�5~4����]�����8�0�5��;��Z���f�:��k����_�èBd� j���\�~�c7��!�b�S���r��(�O��>����iJf;Z�t�V�ў~{r%�/{k�}�*|��d&V��p<�JID�l��}��8��f�.}���>y�t� 9Jl� B�Sl�
>�2�!	|q��ק�ܩ��2��,��uʥD�����Mz�TD�LH.y箷�ڽ�d��r���Q�bхU�>�<�қ�[ׯv���&��W�И�2?�`u���+^�Bp2���u�A�x]թ���U:OR^�.�;!Ah�N��L�u�@��A��?O��6��<��5z�m��"����7N���3vN�2�>�(Z%�r5y�ʏ�s�Rr߃��+]�d������w�n��?OOj5��ޅ�^Yl�.�T������J�y]�`����- 񆾢F�1 �~��A!���;�9��Ѥ�%��&��2?�B��,�_��Lëc��u�3?���a@1~�(�b��tn��2�&Z[�O��,Ͽ;9����K��@C�K���q]�;N�������2���)j {A8�Z�A�HM[MU�Fq�}�b�Ȝ��#�>���m�+86��͇�ݦa]�ʰ��8g`?,.�R���g@�y�ڭ�mt��'\�|+	�X����N�)#�M�%�#�q�:�Mqns�~{,�__n4�JR3���ԹZ�;�j�Ɏ��6 x����cu�m:�7e߭,��1���3��s�Cu�9ll�wiٽ�'���BTp�A|�oó�u���HO9��Ջ�M.g�p<��M��s��=�rh�������)�2_���3�iȩ�c@�Fʭ��VUHF�F���jHD��2�AG�k�f=j؎�� h�]�%o��Gp@����F$^������x�I7���C Nyξ1�9���K�IM֢���m 3�=���^M��x�'�����	��Xᶍ�����<v��O���g�eĢ�GZ2���u����,�^ΗLy�\�Qp1�b�=Ԙۇ�<���F.04�g3��{�|&���� �J�P&�qTS{a���Y�uӤ�K�F@�*p������ꙝ�����ǔ��N��:�)�ף�LQ6`�p	��Ƴ���<�JG�F�WC�S^=
��@ 5�{�%%�1yd��dR����T�NCc��2흶�
��l�sDSW�@l�q��?�
y ���zIؽ"*�W;��_�;�w���._�����M�V��`��{��7�]n�Z99��th��<��ķ��b,.g��ȓ_�
&KUga	E��ɡڑ�3'��Gbƚ�K:}�kŗA�Mx�cPz�}�+g̪�B^D��
�q㑶t1�pF�n���7���*�kq�ZB���4�M��Fe{7����2��)���n��z���+��?�y�'Ns�iEG�5t��A\ٖ�<��È��A;��7O�����Cd��"�*��q��긓�f�/Y>��ԍ��k�6�gՠ>���L �d�Q�O��J�D*��C#����:g�ͪ�x*^j�T �1����^�񻄹7ݕbf��5_~�@�J��ߢ����[���i�qK��U`V�.i��r�7�7v4�s�����qE=���Tڒ�i�(����M7����v���@��]��V+`��P�CaG�U	�!q�e����������h�Ò�V_��JB���E��E��/SA�Ɖ!"�K#~.Yhjhb��n�P֋�ջ0�����R�|G<��r���G׮��08�Q��W�}�;�+��I���,���j�z�2���dZ�DYʈ�qdҁ��O�>���I�):��~ʘx`R�gr��ή$���L���У]��LXu�$z�M��bH|DX)��Tx%���#N�f�����5�`���m	�,ɚ��#P՗�� ����
�c�6d���ah,vw��{Pxhl�n3�[�og�=��m�7�8�K��*��+��_��4Q_{��e�P�n ���IZ��c�k�|���.��{���V��d3��X��7�6���2%���T��6i�A�س����,|��ۍ�`�x-`��A"�A;�D*8\�[����cJ2��Qwn�'t6�4�%b�/�R{a΂*T?��D�,��Hy�眱�j����=�C�fL���s��.7D�Owj� �iK����z����_:{��˗n�� �-�����+Ǫ��� l�$��t�e�8E��CRʋq?�?��6�Uu'�cG���mݒqj��Q�O}�A�HWqF���w>«�Z��t�į�̕>h����U����$�{�����F����DJŞ��}�V�W��w;+XАz+����ʫ���� ��Qt�Ϳ �ggM�<*`����t�Z�k������h�
Ƽ�JL���0]�����O�?�N�ߴ^������� Ct�o�Z]�L��S]��8�񐵺����%^�k�p$��Ĩ7�ע���.#���N�����a�Oj��n�F�W���W�N=����}���R�_ِ��-K+����9��tB@��x�Ʃ,��?	�ϑ���d�J.��u�)�dR�%�(L?j�]r0dj̴J��C�%�}؆���Z�����fҕH�����#1�)�5�v�8�������T�t�������o���{�yE��)���g?��(��Sˮ�)�.c{����e��Ɠc6r�q|tZ���`� �5f573/�(_PJ�x�,�y�T����Ƕr/]Z���Ӡ�<�1�oVj2��-���=���d��X�(���
L�d�m��敚�!�۵veI93�%��x�ѷI���G������a�T�Jd�Q�b-� ��5҅1Mk�l2D�L�I���b�/f�vm ѓ#���o�㙚0N�����#��
�Y[
�*;�E�{����?�������&�l����5����i���B�u�ԑيm�q��j͇S+�� ���3'<`�u%�<����yU4��(;��1����7����x4�-uO��a�?n�8c�����	�"\)�H\#&�߰������(�>Ǌ��;$�S�؀E�&�O�4���fǵ�[9�����8�N �֨5E��S����c2�����o߮9��̾�J��|WJ�8�ӄ:Մ+ _���sO���Yq��4Aʅ�`�<������i�¸��k�D�`8I�W�l�Zw�t0pip���=B�q����%�[���f��[7���9t�o�e?2�&��_���v0KI��;�g�ŝ�,���"z��)�&�M���*6��8+r�]��_�:q/��*0��ivm�#��O��������U*w"sf�{�Y�qΓ*3��1�}{���rY��C��d/�pϢ@Bi��ŔS�n��,SG�rK<���ˡ�h�&�Y��a.����0М5Ҍ�-u΅�rF�-�|�
�E%����d?r�<��	�s~ �m�2��AroS-^����䨛PF���ԛ͂u�#"5Z����@K�*t�������-��!`�j1l����<�~�`�udlbU#��P*�m@��-�&���@з���]��\JN�=�2��:�BQ�����Fv�c �j�gg��e�����+�V�W���j���p��G����&7��Ƶpc����xR4�Mn
;�,�'d��ġ����<���&�̀��#�pݫ�
4�(x�@A2v��h��o�`=��Ij+�� 6.�=�4�����'Y��"�߾����1&��z��١���c5�����c��uI��y��cE��(zcj3����7�47&����i���>�	���V���B��[��=!`�G ~��F���[L1�)w�Q���o*F,}���b����j�imt��,WHd6!��B�8X� �$,�	S�H@G���z�!-{�&�>a�Y&6��(c���-ԭ*NP<�`q<��{���q'�޳(�[��)4��B��E��I�A�Ő�-�syI�"��E��k�8�R3�6��pyl(:�{��],���ƨ���9%�~E��a�U$b�M����]�Đ6ay��B^�(T�>�R�ES�>��TA�.�w�o�
�nҶѭ?@O��S��Koƥ���z֡'�%�a��xz���l>߫oc�	s&�:��H��z=��7��!,¢�1���wFu���y�!K�(sȽ�QC8���s�1�L�?B�6*
��Yz]k�p��]鵬^�����t��'Kw�ʛ�ӖS���}G\q�c�&�k�W���eԅ�jg<��]oA���
Ö�y����Z�<�T�Ŋ9)��J�w��䒨i�����9��A�y�����'�S��9����%�-7�j�ϑo���������DQV�aŷ��S#��o^�{�(���>LI4v&4��C�2��\*���I�¥� ����byN��Q���	Jb���FW<�>ig�.x����W�k�ه��Z�fC�OY4����Ȧ���@^?��5c�q9o��C���s�ٻUa�n7�@�wI���G6�1�%C�Y}���j�d)�-�D���O�"��$I&�����b�!b�����UP�XX3O��]�>���f�֫l��N~e���L#�҄����"b�i���	!����uN�H����)��xa�&�%���te8Z-ME�sr�fͮITqx<���P���2lN
Ee�#+�r�m�GZ�8eZ<E�f��x(9 �92Jx���Qk(X��=���4�B$�DVP�y���V\p�_j\�j���_�k��±4&�{עb�BS������B�*�t��qXN^-�����J�q笫T\Ρ�����=�7�or� �?$y:�]������j�N4�)W%��l$
�Oç�[4�5>�o����
d��ʄ��y�! �K��������K�\�vL*����=`q�������"O^ #}�l�E�Gw����I|""O��79� �d��Z���ϫ�qn�G�9���bKjMi���#@\���`�bm�LU��Z�1iyf+̃��j�K537W9�$?�3���=x��J<)��NX9HGUISA�2��=΀���Z��cDDN����ᆺR���M~�8��c0D �X�!��d�ev0�����3y�
T�q@2�H�I0P��y�Ԥ1j�9����*B*-�`@0�G&?i���b��bn�tU6������غ8�~"�K��<:�h���C�z���'O(zu�l��;����o���{\)im��) y��t.)\��/���=��D���4�eS+.d霶c�
T.�}�ݭ�_År��WK�,�PM����ݦ��~�";�d�1���\do|���l�08g�PZ̿K�9
����\m���伹} ���y f��[;ɓ\v�D3r�p�\H���&/���6�B�(]��҇u��FbW����B͇?�#����x�-*I�� f;����%�iG�}���]���Zfƽa��Tɾ��# �)&���/��~)��3C�C�4=g�ӼX��w���[�2�߰��ɽ$�;s#b��ڔ�{k&u��Ko`wh�|��mŶ��q�v�1��>v��E��~���KP���`mTl��ʱݣ��d#gq�����w��]�T7�zb�8H�6���+�T�|ظu�Fw�3�}�#��X�ݰ��,��Vm^�]f����UG�n�B�5�ih8)��-�$J����f���8|�-�������P�կ�|p�r>��x*(kWmbS��6m�HR�0���H�A��S)��eGBѧ��7���O�lq'�ӥy��䝞�tpUi�Uը߰Fs��/)����H�ȝ��H�QFP��7�3�N�#�6�6���������&U�G,D�Tqn�ɦy���D�\���cAы[LS+�'��kNۑc��	d_Hmu��d�5��3a�ӹ�տLr��zD"��ϗy�ǲ�1�쑽d��pV�`A�o���\�s�:JI�οޞkr�\�x��
LA�R^�Q�'pX) ���N5|W9��E��}��VY_��p���+��hx-\��4_�HgX��^��9�eQ����,���йA,�K�޼\_� �;\8�]�6k�;���P���W�5�H�X욡�4��Ն2&� SK��W�<b4�hFJ�/�ȷ�E��ZZ"4����=��-u��.�qz�a�]����ə}PAα��t>�dz��:;�cH�%7�4���Z��:�����'���s�#���1bn�b.�z�Q;,�\���opʐ@��\L�_�q�)��6w����?��`8J	�����l\u���C�p� �ϰE��u5,z�_&1d8��c��S��P���pD暑I�VN�9�WzJ2о$�i�	o�#s��8?$�)-�*��{� �Q�5�cS�"��;=H(��tT��t���wȵ�iuФn�ͅ�OaЄ��Nr��䠬����b���3l/�����C�ԴĲ��p�&z��޵����Ur/���B����'��s5&;�*��*�$��V[,��G��x�қ��$&v���N}���6t٨�w>�mF\��x��&8����6�G{�/�ɼ��F@'T��6 ��%��5�U.�G�����.�g�
&��C�/;�>U���n4?%�$��Ry��k�J�5�?�0�hnT\*F2�"��ߩ#�kX�o(����u��f��]���D�/�c(��Fw#T���ѡ��C�M:���3�:㺯�����3��^��Z�/�%�qC���zh�	ZAG���((��8i��(���qß����7�Z��!� ��9�e�WA��(W��k!��~�>�,q+�5Q/� x� yL5k�cR�J�l��P�U2���W����*ie~l��}n��-��]v=���!����By�d�˷ {�K>�3h���ᕈb�἗�#x�Gڣ����޵�$ \G�4l��+ȤA4�I�=�\�}�4��u�31�	���dЏ�L��I�I�a�+��'�v����j�/@�ɜ<��jՄVr��E��+�3��)1����	4��ў$�T\��h�v�N���0A�uS��۷OܻCo�J��q��ټ!�Ju��N�r�&otq�3�_6��G�t�I�7�4��M�o�z��JԦ��� J�C�J&9�;'m�����qv^�ɯ���z�y��
����:̱J:��8_h�O1��7!�^h���h+��ۜ�wjD3��r�"������G�U���2^���@֓�GN��Y��>�0��ɨ&w
�8����N�۴(�ً�g�{����$�H��r�/o�v�g~�}�i�Cc7�H�sw-�F�9\�9at-c"�**��-���?-_�RL����ǘe�^�x.��x�Ձ���\�zGi0��w���-ԃ�����ѷS� .��!4nI`������(�a�!k�A�v�#��=���2P�-�Q�/ �r�`P�d������E��V�R���6��P�ܸo��=�ƹ��*p�D��
Y;���������$#04ȔZw�sxW}:{�(BC:�p �+N��v�;�Hf�6�U<ܠ��8�&�'�����E<��YU�?��A���Y���a3�&��?�y9�/���LA�+�p�	���j:�F�!�3�uKI$}݊�e���U8B�mЇ�L�r7�kr[����i��r�t��W9�����A�mU�UWEa*���v�X��૓VX��
b����Z���}iޫ
����/I��d����N��%��^��G{���y͟���`��=;J�[j�!El��I�ތ��z$O�'���x&ǻ�C�ۗm����0���y����KY	�7�  ����,k�OEB]\]'�r�H���.����p����ʿ�*8WBN��dt�,���G�g�	3P�>y�{(`1%��nu�b�TU.'E1K�|\:�M ��l�M�X�&�hn�XɁi��K�)�`eI/�sY�刃�v5�
,�3��^�=�s;5��
uzLl�i��C��Byo��%�Rۿ"�bt㯍�Ǖ��]���� ���p4Q���b�(na��3S�J=p�B�?0��m�IF���γo�G��(�� %�}�Pn�%��z��@ҴM��gR��6�7������w=)ϑ7-�ٴoS�<8c@�6S �[	�=�kmU܈xt1���JzQ�d=V>��[!M���#��?�	ʐe=>��-��:�ԢQ�����Z#cd�v���T9�ſF����K�EgJ�L5?��gH�w�����@�w����ۏ�;�������7|>Y<aQ��:�����[�0���@�դ05M[iY!t��{�����Z
���9Hs�	jafl@e;�ej�ڑܽL�T7�z#�7ד?я��5�D��{N�ک�p%'����2���|�)�09��p�_���jf^��<�$�����%³�����u�M���8,����r��f	laMp��U�!z�S�l�,P��G�L��3�d��[h٠�\ޡc���4G�{��7W�w��$�*����aÏ�0�Ď���C���o|�-q�ט���}h�� ���WJl�$E���AՈvj��FibhCZ��V�))�u�D͜9`DX+� &�B�<4O4˰��B�Ԏ���
z���t��#�A%�%�h+
��K@4=gh�Q�%���oX�n���&X�z�S��ў��|��I#p�]��,�#$�jh���Tpof�ysZ�9��@� :;A=��E����)/y�D˥ws%��nǂ��;1�v�J��-e9��C�{�Zo|��j����1�h 7�����q�,[����!��ڪ��86�W�ͭ\K�b����(�-�i�y��9���\a\�������)���{�$�O�'5�\�Q� e��Iz#���j�ЁB�-_���Z�D�"e���ܺݩJ�R��VهT�J��(���d�C��\C����Q�JyC�q���xd�Q8]O:�F���pe�?C�MT�m��7	��s��N�H�c��>��#�T :I
wǰAA�`K�\�F�h{�V$/�9�jU�c�w���(M���-�'O�h1LM������Q�&uN~�h|Jl(~��@c�ͷ�}��HШ{e��\����U�H��j�%?=�m�ap��Vo�j�mcH/W�׏דh��	���?~4��u����d��D�V��H�h_.�3	����A�����&��,�[�ZJ��j�WN�����'�2Ͱ�Gk�I��2���GuC��<��nw�Fo�)
��M$ަ�<ª_��@�-�GzQߒR������w3�q�]R,8-d,��+p����t�c_���Ԗ�=_�uU�هy���Zlgj�b58��-%p�#�d��|�����wq�#H�Q	�4�w����y>��fP�J$������g�C/ɷkE�cK7�?@<�R���(~���,V?r��/v�ZyM�q�+�^8�f��/U��{�7c����V?4��Ԥ�E�Z�y�yV,�����a~��P^���E<��������b�t S�F��j�&�@��s���+���c[v���ɬ��f��V��Ե�t>~���xe �^>���H�	32���$J[�q@#�u!�{�r_5-R��t�L��J��1�TV�}h\U�O_ϩ���ò2h0�l�J*����;b��E*F�7y�S׭}<��=P����qsQ/^��ڱ���j@&�^��ѪLO�� ����Z�����u�,#�-������[g����#����e��2X�{�pS��z[�G3F��D+�d~d'�h5.��������j\i��1%G��{5�DX�Z//�����u���/���$�x\ ]p?�Rf+-�(��v���m2��2��a�U�m��wض�U׉��J��o/c��A�%.�2�X������f�5��\��(� ����tZHd)p�׻r�]%U�1�Tpz9�X\9��UԬ�؈XEm�E�N�?#��a�F��d|7ϵ�G����+�T�9�Kjd����Դ���a������l��'dS��ڢ8,�@�=-9���,�K��1X%1O}M3s�($���7Acv]�%ʦ��W�v`�K;w����ȔL8�5���PX����)���Wv1:϶�V���C?W�%����R�m�3�q|��0v&��N���H���&���:��ڐ�Buɷ�K>'��]�=�Fe�����'|'p�3Pߺc����jq�&�;N>*8��O��� *qk�9N�0(v��I�&/�tY�!z%��)t�)ڻ�>��p�L�$���pwk�@�aF����U1����ś�G�Ӄ���y��bj��+N�f&~�0��u����/6%��X'3g��hE�õ	b,(KdYp�J��1�3�^�'��E�Ӆr_�rCg��<�J�
P�5�<�&vf��7���q�Wu@�ͥ�zz�؊�1�l���5��ca]<{@s;cU,���;��M��3oa]v!�(''ԷM�F�ĭ4��ڡ���Z9�`�ͻ���EM�ϋa:�q|w7�ٚ��f�R�1�
U�w�*�����5�_l�6������޸�oba�g��]�k�� �슀 �AXF5	Չ�B����0��3���
E��Y�X_j)���L�ǳ���Īɶ�-�7	}ͻ2"���.�y!zs�o	��Ac�^��dL�R�'�n%|�
�S���:I���rM2����6���Q�R_0_L(��nu�,$N�(�('�y�EY���X[�$u?�3G(6 ��F�ƱW��d����Υw!�_┮Q���/�����%�ǎ�:�y$ !��޿��?0��yMCx��Wa%^ey�͸XX���U����,�7�E��Gq�`�?�B�W��r;�m7O�;��S����Ε6V��8Hm��;��Cs��lf� ��2��J��)���Y=��t2m�zo��H7�7�	�M���d��u2�9�����h�|�j�EJf��y������(�#��wz8k8#L*d��(����]�ͩrEk���Y�o��qI�������'7 _Ѷ��ӓ�ܸ�5e�>�q�!q����e��)�ףi��A����{{æ��5�����DT�����دd�T��8 }�L���,�4�+����:��0BW�˽��,�?�}� �]�/�V@�̰��?��g#�e޻�K�X�7 !z�A"��������g��/S���9�o�[a=R�@����5�5��sP*��L+Q�E��{A�f�7h�X��ms��s�]eN�,cs���`F��\�L�ij��t�cW�Uӌ�;�/�`���k{� 쵆
��M�a�|�B�F}g#���d�A�9����R����t���V�x���z�gG\�z��B�#�͓�V�P_-7�� ��cXa������D��h���x��{�f�)ӔA��?81
�L�krۄd��f�$��9����.��<FcG0S_]3���d�-�~�"��g�nz�/��U7�Y8���]�~I;��0�5	��ۤ@9��K��;ə2ׂ�]�ӜP��{�-D:�:����C(e<E�>���7e��Gxq�	nh��]��^��,�����8H[N��
Q��D�g�@��}��
J�p��E"�ź��Itz�G�͐�:�u ��œ�A��q�`\X�w�Wv��Wz\
O��|_rC��j�ut����̋ٜwK�#Ey�OP��"h��P�융�RlS����L%���ާ9��#<8&�2��hTp�HM{�y/Ĕ��!�HcXlWi�8�}�T�L����0���h:�pm�t^�j9�IU6sV�	�9���,��U����O�[�,3c�,my�'�1�f)�5U���\���^�Ψ��`�W�
�
(T���B�였ds]a+�L�-�j�k�g�����q[m�q�qaI�Kiѐ�Q�ͼڢ��[{�����*<���T��}Y��m�-�}ۧ���-�c��O7�V���(�P<�5��K���R�܏?���h���\=:����}l|�E�����z��<f~>Uۼ�B?���!��o����X�]��:����՛���h`!����%::7*P���vj����(��Ӽ�䐩>0<�$ui���s�9w�=�QyN�	���V~�ۦ�ŗS��#:��f�ڛ�]���K�:>��pp���7ƈ@�#x4}���B���lJ��X�7��F�
V�	S(ѳu�Ԕ���v8�	�[�ɘ�O,R��L�ǔоD�D8���{��{㿙qw3�.Ԇ3�8�~��A>	Ҥ�R`�,V�Л��>����4B�HSO2��l_���+��`RprS����"x�}�4�bY��a�V�����F&:(��z{��b�AV���16i��Q�b�	��'r� �����gc3S��_[���F��T��l],ݱc�fB}�ʒ���Qh�7�*h�Na��JL��ZȾW������/C�'FؙB2ў%�0o	9�Uu>䦢(`�u��E���X�X���\�H� <RƥC����cȭ(���۹^͞�dձS���p���W���&�;Cp�gmN��QU��J,���7#�"�����.�J��ѷ�q���O?0x��(��~:DyS��<Cl�P������ L�	��O������g}���h*lr����?g��u���8�_�R(ĺC0�FQ��)���?=e���ň��Xc��ўsTF�K(�9f�%����aQ�s�լqM�5�\`�EE���~��w���Ҙ�oi�B2�dU��������f\�~w+m^5�jW�(��5�N����rU��Pi�((���&*�6�LY�E���4�C�|�dS_Y[��3|!6�A>����nGϺ�Ak�
��Ȳy��-�[O�ʲ4k@�it��-���|�ֻ�t�Z0�W�2��5X-Z��o*�:f'�Wu"�q��NꝚ��<s۲�><]�!����#CC���'�z��(�u4k�����EgQT��&�V��PhS��&��?�fE=Kz��X�+?��|��b�_6C�OBijk���U���$e����iv���s�U���#��a;�U�t��x%�ߣ��+R���)�^8�v�Z��ȗ9�[�B��	��ݒ������0};(��;p�ˈ��>�WX���S�MF��W0��p�z�Cu@Ÿ{W<�}>+;�M"j�cms%�2&�y��M^/xt��vgJ���0�W}�c���M�o5#�.a�W��ۚ�W��O�/��9�����$��D��v����XS ;�����j%�1�����^&?��H�jU�����@~�&g��Rݥ2e�}@9��To�"���F|�W�J��Xۼ��Q�ЋtЙ�!���V�7�2�!����q�qMѽ2�l���HŐ�a�-�������&��B��m�TWv��t$��[���C�Q��ӣy*�6K��j)Of+WǠh!����>oxV�h\���%�G�w|��7�H5/<l�p��d�����K6���S==���
�`�kC���\�,���}�T�~>�jr[='ڃ���3�J�r�TQvǈ��}���ol�.�s���Ἰ��Q�pZ�7F�c���� ��3B"g�
���{�%�X�+z�s��<��ϻ4�yw��Y��$�n��K��?�+��E�� �/+]&������ʔ�։@��n�P�-w���7q�@�c$�_'Z�A�;W��#Y,��c�=�����|w��˻S��.�Kb���<������+��J)4�%FZ�4�sP�*��t�;��|"e9�L1F,]� �V����-�/Z��*��@<�h��3d4p�HXrl֗i��ˠe����D�l2�u�ĕ��Zu5��l���s�/�&E>�U�&� �%�I�+ �B�'1���d�W���j;o9r���d��-��|DP+�E�
�)�wM�2�%�h�a�(t��R�ˍO��<���)#F��م���FC#�}��,��+��3���c�h����[��
]ٗFHt�!ׯb�o$�G]ہ�j�;;�p�5@����g!֑�,�\���VMN!E���-�n�w�7��~ٍ
���ku�@2�����`�z&��QR��;�W�0;�u�G���>]�s��l��h�o~Β/�/wR����Й���<2���b|�������Mj!a��T�8Ob��%<��S1ȵ���O9��)J����3���G'�����6<ke��t�9�xq������~��eSn��"����h�XQ�*��4yQ���Q�ld��.�Q�0��b�O:������&�(����LU�e�,��`Ov[`�eC"6V�#t�|3�51~X�g>�lDbA��R��ʐ�̨IT*P��	���S�ET�Hh����e^��Y��R�w�Q�Jy1�7-Y����9VI5WB�����yX��n���e)��)�E�U�P��N���Ӿ4L*���H��i�5��_�[(�!<G��P�$2@�W��o������qꦃ.�&e��������Ȥ��iB��fޑB=<�1�������0K��F5j�����ƹ5�z�_��|@R�6��p3���\)�<֣��b��.=l#x+��
}?�5oދ��'�֮�b�둫UP�LbgE��|	�~�8��U�o_����:����ڌK�@h�82��։^%����U$���P���x{D�}�u*���I�+p�&�����)Y�}��*Y �7����co��X��&�V