-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
V9nLQ6fS6RntpjB03bQR2rdw+3PdM1SAZjuyWB/D99rDKwgubCoV/d9lK9gAcWi1J7sJBbSlvHiz
/3y6dgYXqgi9g6NveW2WUzsHLBKkxHHZ15i2PzkfvsWOdNNZDuBvhZAWFBpBgY3J8t/PqNkffwnz
fNJykckGPni45NVT4jgn/dWXhcGaGWlppaUQhrjB0S3wrRCGh1Ut80brYsmYST1RQ1BqlBPurJme
rrsM2SMYIqbcQEll/PoUgsKqD9GBhplGoaKRbVdpoq73YRUF8Jdh+aYIw8NsNbkUDXJH7gqSzKuI
VaO4CQgT0yyHfEcsNGSyozDUVV6hW6uTBOIloA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37232)
`protect data_block
5mXVVWwxSBH9FSvp+kSxSoRKDOYIAeg5iGEXDaAGPqEN0zjOMN4JFj3AEuob8RcnEIm63UBhww/5
/EXpCHGvSjQO1nNEWsS6EhTuQ6Kub2inS+LueffgPajoLuCyONTcueGL2v+9pQAGbEpPh125LKDH
91odXME6r8Bi7zvRYfZaNNMHG4k3w7IqhjSBT+Z1PyWiOPl4eUSFPmfXMR+rmxEyMiJH7KjaGT7/
IZZbwxKJ17+DF6zrJuvssIijfqyQaB3PcGjHaSRr1ttzrH5gObYQjI+CawIWqxM18k12sWsC4t0S
5HeRJzOQt1+ma8dBu++vvl0otnAXVBGWPPCQzF5ZnmzRrD4TPxfc8AfAQvSH3sorgt0BUo9CKn8F
nIKbB+oUFFJYAKErtQlwH1p61C/WJLG3E4CIvm3Bw+6iyzYeklS9zOraXkoJSgvnXvcDZka/WSRf
P13E9hQqFemXQR8EppB+29b5fY0+AH0xrtaI1Qh905NusQ0+R6Ay5MWtHc1L1TTk3pNQJYPk8SX0
ojb/s82YM+Xeo0ze8GRJzIxl9lKCA9YkeaUg+pg5uWaLPmL6inl2OAALatPqBMdew0VZ2oWtQvWQ
cuYa9Q9yBFE/6T2CLKlCNK5GhstdVnJj79foWhQjWQzd+ozI3jjrPYMpyfB5tHsZjbfy3OWpGVc9
0wkUfo+OMWzsv7r6ZYtmJUP6OnHN1IOwo74V8l4jMrizWXdgA/WUN3I2MI9A10rCkUKjIJy48ABB
fXKZ+oMetfuR5hDEZ9EKIL6ScujVvVPucMiBwnpc+Iuq0G99XENhb3jVijHVVeOaaJFqkj79JOCq
Y5zlzTenWIFFZYF2cyeApoGBYjboZs5hBT1b7J+gABQ83NnQzFB7TFdQgmVYOzYhL90pL4NzypRJ
dyVhLoWv5hgKrzxDdnVrzm4XNc3uv7UwkQSutonVB6mxB3J1JM8QYgb+r7BcxBCL8CFlwG3RAT7q
3KNjwmsKU28G/MCxZ0s4rxtMGc/KVl0sLMRBj5DhD8Wvp+ABA4nva5zsQQ/GGg+4IZ7XgUw+Cc8Y
++VyAF3Wj6PemNxZdcGohUlJDDqSfvzJjFVCRMs6j6L3WZ0+GcPxdnSILtM3jw8j6ScpqY6xVlER
KXevdtVRh4BwwQ5gg3w3iOVqpoZ5weR7DPMSX4OW4sSEWuEmm+/7N8xnly5L8g88gSyutk4R+PG0
2TIPlWSleRhwHFsPkZeWr1cEBuQlUEJSEJDq4zNmmiOzNnXs4+0NznbX+wZNqUxTixIvIQX6sryE
1ImRMZ+Lya7nLu1mzaDJ3+dsr9wBHA3neoCcHkU3ri9ofuqyj8n8nxIPrjNKUNTpR0If1BtU1MLf
a3qM1RIHV4v+W7kz6cIEAwx3ttuNh7xxRrtmkBThRml7+JaW1kRZm5SSNJFfkSsfG9q8Q+pIDR6m
bA6uXbA2nO6xBwk5ciOwNc1eifsiCrSlIo+aeXs/jw6Y8tPCUJ266Ylrumj764MGJktvC8z3y7nG
3IwVxz9QPAWR59c59ZvVfepgaS976gKYuFy7m0hvHTgztFk0NJpOJG5Rzn3ErPYROcu5PqW+kcl4
b7soe8u2+uh+P1cUnU28kq2ga04/jJAO2wGJO2zZbsV0ruRXJswEGwTi6JUlszKbSy9eF9Z/Hnv6
Ckg4oirxGTJOlVHG0gQqkG3lf38faPq3qMrW+1ULZSUqXKQolz/EWtSXMwOdW+yHZl0oCEKZgJOD
JIyTAXt/6dsH0L5HQ/eCW7aeD00gdvKmjb2gCisD1DItnCrz2jgOtuezb+nmasXyrGB5P9YZ2Jm5
lXd0cEc5SHfPTyabhg31SUpanZyADbDNDFQCeekB+LOlfkebYArCQlBuqhmtaDa/7oaNMoNMDgmT
oAz9Rs/D9gMzcxK8QrALJsQbPgQtNoepk38jz7Z2pLOEAVnE7AnH7qllysX6us5CXQJSu1IDW8JU
/pQVBL4K1u3TkuvNrm+Ki28OeZRNBbgp7jowN/2ZHgDoTL4Fe6hLl1Crt3SGLhRVBxhRi/c+UMQ4
+Qz7XvbgXtydnpT+u8WhwwBCVt6D9rhuOn2A+KVddn+7aeo5Vpu3D/c3/Sh4fDRUNwpQDMoQGUst
hVTvgO/fly0j8cLmZj+4u6tIXgYYuoHlD7AtQOqGMFx0NNkKfHbEV771mNoETjnNLjanmNcr2m77
rqDE3xG0W5GFsVWFBJrM75GlxcmXTYUs8C/Q5Z7X2LhOtiFEXRGh38PWMen+YLYkSAfl+YWxwKCZ
OXuvMvZelZvaxm6tbQkE8Urjl5V69hOe15i1zW4ueakbYJF9gl4j/3TlBZTVeLx4a8xKnnrFkzlK
uSfIQrPMxu9SuGTUU3ttJXr4ugeUld15RY7RE5akZ724z8HJPPBh7bk8ZgFKdL0BcaVvxYylHmKw
Hx7CqEAW7aPO7EXe8lH10zticoAp8AB1gJ6uj76iMMCZuvgNo1ASjO7PHKco7Oi7+O3rto2pYYKR
1lYe9fQRRCe66RIrUoS50fkGfqlbC6a/JmNf41jFg4pBIuEcBuKs0am8k/batgl4iUCOSwOZNwU+
pzutgKIOFYQRucoGGegvYCvxc74CRg/5PTv+bN2s4taxQ0VEIGuQmXFJU4lrGb0pj9wWGVE+Yw4a
T38EQCRwIGXi+7CiFgGs5z0PAsB9HzSn/5RPfXnwa+JGdaCyuRx7EX56H82zT7XVRrFTxnK+6TjL
6sBYnLvsCy9j1Q/ZRo9pycHtxG6jT1CsaL0jdmaRNNJ+1i9JFl4EDmFFQCxai6GUk2MnPAUtNUOQ
9S3i4mwoQp4m55MSlDHPsVHDYSUOC0PMNER0yCyCqcRF9jgAjS654XhJn6e4J9QcJY859LDY9APK
eF2kJLkk2n/DrsAFb/cFrhD4B8y0GfVmkugpVsUR04P7/EZsBNksjYmkA4S9WXLmn3SIfOy5yqEc
Z9c+osp1ajjcAFq6s2vU92uLtf1Rrwz3inRGx4nkj4SDAkX47KybYx/F586bENG9XNFbwHU3KZPW
0eycS4s+P1zir+QmGoT3MQl+Yk06uYZa677MQRcujUR9BUAhBQlX0W+EDWXAeh0vCK3WbU3ZEbNj
ug2nWZqpTNRNIH/R+crlt1/8y9ztxEzSQxsdTX41wZYRyqNiL+Fu6dH1Fe5BY415eCz0rc4MpJ3a
gXyjdZcrXwFFWFE9hDB/NG1ZBwVHnWfCVw4/aJy8ahBRVn6SZFseN8RctEdUp25lqV4s/MAuoriO
4o8olIIQi3lgydt+Byy9Sf6Ncrsbos/4gIInSrLXuSoHucoXIsFUgLxjE1X5cZJKIC63pgGO1RUs
2uuRfiGkzbKqx+Z/Tmzm6srMd4ixt7jkqwV9LyhAhxSqp8Xv5RhgOVTCNFT9aSsUgTKpg0fAREsi
GhKFTFS6eIaKr45xlyIVFl7V0lRo2AyEu2OrCZIjR0dMmO7EekxEbtSsnQVn4bWSQoArMB/ev0bW
0K8Exxpn+VzkeL5lbhvX0ZVpxte/lQZ/BI8xUh2pVJPr/HvsPPkrya67Ed0qQhQYmzsdbGHSsI3e
KiI+emNFQ99b8QXZo5S90hvJz6zzvDggI3anx5HP51PQoOatzsX7sciq93t28ArJwOFHaE6wxgNm
9PgMLV56zGsc9B0zzh9iTPKMx3YwAvI9mvQC8D2hNz85bIrWgf6RvLIvcFOGQuLg7BAdtT2JlGpf
5KwfYTlPNWIlVlEiLzcXvbrmnEU0xYZXNWt/nl6kFWWW3/UHElJRYFOIOhcY2nWn5CVGGSPbE/z2
E/qK2nVU9ayhFz6wd+L/182dxZlUiBMrBrjajWhRgCkXWlwZaKTYz99j+BMa7VNYlfLFx8iQ2IuD
n7OXnBg7IfElm+D06jkqeZBBh5vX+qdl2/rDsrdOY32V+WJ+U8C8PzPFQJ/ekAczsb8u/bKxB+UV
evfmbvPjrNYYitFDarxr52gX7HhEgXufpAYGgdrgrUIOgVwh7IGDnuXjiCOIuFyh/stKIpy7Vbmy
JeQqPhee7B6vu7oqsG3lLVyXtoAa5v4CtwMKispy/9nVO7TBk1/n4QM8mvqVezUIPQvEKvvlB/QY
d+19cV2sL0nC4swuS2F7WKwNHuo4s26fwWHdxiuEHqnn6MGRutuscnKzvpqcK9mDQurK1ymzMmA1
S4trlu3Y/kKVH30fZKIeJaVpCWWQM4DWpH3XxMcYH2ccBzZrLCTXdFGfPb51hyBxTcxsE4M1WmRL
gUvNRUO1T8uVCt6gQZISX+uKgPqMlZOLggRJ/hEx23YXXNBL2PT3SFTnTyDFrjLOo8Z3cBcYueM5
q8iykEUeO6R5QTHtf9DC0cItE1TCAwsZIJ4khju4PYyDRCJFGFSCOGJJSkyzCgAb5IBzOGZYO6Xn
DktbhYnopC7R+/XzG2nPuZO/7fSwcQIojgNgkcuYHDxWUT1Bb36FdcMBPx6meViu0WaQ1qGwfylx
YpVnHHWkJmgrIOnezEx32XYlj/10PQw6EHM4LbrxbB+wdzYzBKvlv4Er0YylRyaPeji9mUdoLnuo
2XngoPXIpGIyFkhiIoMDlet2maSAwF8gZ/6GaYye3PdyDQWSkoKU4HLbIhHugNy47dIrWxNz4oNO
Tnyj0d4tn6Ooph0X1rkO4XWXYe+R9kMJkCPp2mJm8FobGUkgv9jbOP4xK5NIi5KzY+IfKxkDaumn
p/I80e03omotNbMx5+E6quKra5pqQ5fElZb6w0t9slzLi1bCsovUoQ2cxtoWVFRSJ+WZtscFmE9Q
2rW0o7YgUu7MCbPl+hgf4nFxhNQo+Ir1rBXfPXS2VfehetzZc45oF5QHtKUZVMI6ZpEknyHuHLl1
iaLW/vJ2achvFkmHTbfvEbb/gjvyAizzXc9Du0Xr3MuUtpJnQ25wpBzR8lDEpTarbAkjbUQ0gIPu
WcoNoSu3TsNZT1UUcDzlVS8mgWlXYOB/ByHR4m3LKz5puL78OtBHfTlbIHoIWZ1conVawxHP5g4y
S/AqWio/ju8ncH9/V6whcx7YERx/Hwk3dSZopbXwFTozbXOA9lZQOFFU6U1MYxcRcyGsuslSqzQl
+m6wuQq+F7di2BFfxBlsn7jWkjCThqF/A78BFPP8BS2xehWdAUMz0y2ku8GGM/mHCaWNaHZWQArm
7gXU+ZjhpwbQ7oZJDR0QfZdJM/Ib9d599oSIS0VsFiMLBvk/ctdyVfaGsFb+xeIIQs5mz5px8eTz
wFZHL2nKThEqCZF7bDsueipgnwoSRWqrQFvaPcez64nTFI4Uw9ObuGCoPriqNSP86ubzPxcWAxoO
WAwFnwQrCeCpxRUwPfHHjIMmUra4wNQLG7GccCUuaxHbkNQVxIjpGUlnEdqp5sz1trlWX3WdPBpY
40WS8K/zUEBb/nFftM5fQdZhEkzAZ84Lqjc28Wa6uS50pGWnLEDY/OyCWbpMCqA/a9a14sGRjFVJ
Lw8RD3/iLljnX/0jC2CDaQGDwNoXrPrDUhqFKSUBEOk164WDrozC8Svcy5t8h8fOJaakzZCFNxhN
0jobyMhemOi19VxQOVt3JrYBUdMgTiMNWTvr1pfjdT4nd1qR2F7jQZIt4O4eJ5YAOG0r3akUTb5Y
NIj69vMagsligwiBze/da1AMbZf/YLc93XtDP1zo8KJchgUXqHO7ZEBDeVRny+RmKQ+XKm1YkHSx
7w7zTF5VzisMQ77a+GX1S9Snh6hCIVmDRlW7MHwxa0URZuvwt5Vn7L5SjQzh1zirQX68dOsperET
OxU5aYZDf0Piw9DvBbby7c/sklAjCx3d+EyezHR75UrGonfssud8iweccVDOpdX7apl4j1QEpA3p
W6k2O1Q8kYm1n8EW3updvuJ3QnSJI/yBkdzFOQQB9LwtTjGJ3CN2ipPxhgYdb2mW49frioaQNsGZ
xOGsDbnYu+OHNxKx6aFZLe9OOoHjuxpUPLjEwcUHmYZe8MxA+c5p6qZA0aLWvjgDk7iPr4lQXMCc
CBul9Iy3WOMpgE4XZCF45R+jQWT5JeaQDBkK4Xlx0NQWhjgGW0APGqexRGeshM2MRl7v6sWZxg12
N5mirRT7RpjczPRJ1E6zltGasHmqUWD+c2InEuVetiob85aoBaCr5Xfd6BI1IiAGBgCw5xYibMX8
HgslK2PpKjo/64jCpsLUHkb5zxDEij6uL8T8vYkgNbCkpewkhGPYKJK1bCgUH9m9zVB2Km9NXvd/
qcZrk1kx+kDNAleQGfxzwWav41qdwVolDyRprWr5qUZKEpMmJdrc2wDDGWvxXHcN2KGv34gsLQNF
vnLPnxfb30WJ3nd6AWnq95OaWN0CoHdCUxkXtVaUzFLqztnyNgH4c7530V5tEKvRu2MCNCaA5Tln
uE8HjgA1EVsqoC1cfR7cjH5srSzlB/yqoKexRIvRmaDRiEKd4Zply3uyTNuwYOnOLWn6whDZMjtd
zbkjCO2vvoNM1t+KVYBOSmgpBAgo3j13UzsdorptOQrTI5ZFY49jKYHJaT290WNCJeUjRGytEUEY
+yiRJIJ2SiPE8cIx9SQ9gAkGrDRTgXU8gSUBcwBO3uKONbNCQGPnRmZu+n7HSOKHXFuSZcOKWY33
aQwwe0uGbUKxoJtH7nBJ5rxst9EBWaa9yBbvY+Y2yUT4T82Bn90ClKyLAYs7ByBXvLIYIdMAPwRV
SVOPXD00h04V0pT7B5XOK5G3g9+6GJNsgH8TJFKmJntZHt69Od9w9DnnLYRCLv0nkL8guF7LbO+t
+HJQQZ59oRR1D19wmQ53Ktak1aHcIgbNHLAuI9NWPh0gz5S03PORTOwxUNw0j7wbrU3Fk3jUsrf3
GT9P5o8OPjkCFDlOT+qw+SopawYyJBubj687KhyHri8WmlsVlsSQhwocuErsjPZc67qAk+pJ7T1P
+mOd+lsuL+KCu7ustk37ucMDjeqqzW00CywGdZ4YPfNDo6E18unJ5m2v46hFt/y9MOuLxBJo9Qrp
GhTxKjxgQT/g4J+Hu14EChO2DmqNWEVNfsCmlvkZz5egGobgFKRorBP9wHLdMVqIwMpye0ztPxWq
m/+pVcbcijs6m4vBygH5UDXv2qvBVlVz1vKyQMmM/4F8WIJVoovcnBKAxDUqyfVGGAbVdUyOFUMf
OMLI4No5NJdzTNp1nGbUgRPwcuVWBY3leLEc1mFeD7b8b8d8sVvfanXmPevRYXTxNqmnnj0C1LXk
Mx4/GQuw0UtiuyF144Eg/O5aF86aKfTSPvRXOTIvNPdhEA6rSQbOSC0Ozfow9WgeeVnKr1DQzrLR
3NLTblk61EYBFkve6Bxs72DizZEj93RvD1qRDv0DplZOrhzf0KR2kQMb2YODbWfp8Kgppl0JZ7qL
XdKptrlQ2Ktya7GivO5YVU2SzGBQqkfIJeiaWBC0UIOIfBhdltcKxiZqzLUnDbzMlU44oZoImoWo
7tyZcEWZccLGEdt02eLmFLA0ITSRqYFmxSIFOT8Enp+0wjuUpZ60VVPufTzfwd0yZAUcVsQqWuyj
jhmo3r+YeU1oHJNmfgI/j9IpeSFHr25qDS88oMuA8vxKDPUsul0Ms+H7Y2YuS/h0JbozP0zdRKcW
5k8E1hrFpJO8/yBaiYRymyv9SZB+NnXF6IwFRivfCqCYeywJYZTIWER9pfuGwHCoGtjRwKu6dY9m
iVAqbD/JEF6LA1u9xu+Ps5qm0ha6ifG+8Arivwf2RqqyxQ08UeXW/xPxmrYUfyp/jzuime4gjhBi
mrfUA7Nt7KHG3M/5min/Z7R8z20Yi8OvijgJw+SykfDHFMUIcVBbp2HdafYzQz6b3YqJ6MXUv5gE
vGxi+ImtsSsaeWlxEDf9Fh4HujaT207/etNXBcm59JH3wY2P9fZ1p6+QtwUlBWkp1w0QWCxQur46
BxM5jUmuiQPPKDJgO8PJVmkMIckO8SjmGx9gnTeoBb4FU2zZDth+f01dQJbB0t3m+tVs6XjixrPp
Z2N4ItT0UzjmwY3kjjOkERybFr7ctdYBHnBG0EV+8Iy5XBvpzF7lQkjyvziNQVklMtJ02EcHf+oH
vxHI2Jjy9DDjGKiMKt8wY2kTtbpIAoWt2xn40wXwEgHPPaPGgqtVZMN7N3IOfcbnDT+IqB2QZMzV
EpmWUO1p35C7OBt26xT9IIoBaLlRl2N+2PqE0WlLdSLOFFRA5IfiGJOrRSwjr6hHLFBqE8qr/4rD
nuLuksVwUQ231hJayPsq/gH0wTa47EeigC0JeQyAhqb/2dx+u1fYEX38FRHakrhE3+ORAToE+3Z6
g8SQ5h4WC2AkQ7CW+2ihZW7oFWhOpSVDdl70EnLyZ12T3BYaNFPulGs1UbcToswh38rr5aKv3wvs
YZrF01Y09I/Mr46Gv+NeiwZ/LF5hRy0jcsemG7bFt1a0SyLsF9jZCwdE7/TCnavy7KLbnFa4Igsq
PqrkmHiB4JcARwZwGu4hAxfchcElSGi/D4cHLmucEbK+eeXtGV1RN1xrmAnyypJJ5cUyuNCSGzJB
sQEe4XwkC5RjXbbgEYOwouQsxuA/qF7TKoJOEyDc/YfM5FhvkZvzevj80M1lFK0/nGvZWj/30dzf
7H6SqPtl0lIilrqNt/btiD4JMpodqIEpK2dDJqskGoR6BW11JzcmriGu9x4sYgMx8vYj3aXWp3fz
jbGsxnCrADDKRbz3O77UNb0pvnSUwKBFXTNNbSTzNW+d3RW8oGpAiUpl0LTBMU3L+2+XSxj4aCPo
Yi+ocd/EmIpU28QtBRHXFISyIc5lpUNHDJolrhVolkPqEfRcml6OaZqleBswz12pGeyv0y54b+U+
v3OLS8TOQUuKbNgy5m3e3piNB3SaSuwik/1M4WfPS/viyUjnhHkg9IU++WaYrwFn1LM90OJHpYlX
ljvkFvE8KvIr4XVVTYRUf4ulb1SUBLzfGZ0bAnXp1tXOJ32zhn0c1/Ib2SIbPMBMDaK32ZcbL1WT
I+jU3sruHHzmMCKNxPK9kKJ8oiS8Prm3DBg6adp8y4wOaoGYZH7qZ6xO47p5xjBEHDWKu99td+ZM
k8iWmXMWkUOhw0Vqaol/HT1dSzwwmaEOxwnwlZzh0MJ0PG9Y5rrVnDDi1j6W12pTlW7eMy3b/KpP
17pFQ7ukWRjCwwczaha5UfG5agqYRo7EXOrrMCz2VTjjQPyJTB9Ympf1Fvjy9SWInvRfHGFbjPAJ
PxEeOkjIIXfX+Nz0nuiMyRgvCNpSmJIBFknj9ZTZpPfblNIx/ogS6hhQdV2HVfXDEy7siUBcKVZR
fB39dyZLnotIeo6SrkHx51c8gRtorsq+NKKrA1csCRAUuCXsu/cPJtVgy9Y+SlTbyDiIwCtuE9Xd
kpaX5d7Z9e5FmN3cJvhhBKzUw6HajDOXYVBNEh31F+iXrWtRNT/oE/4oodX4yGLOJGoR6M045gq7
32AaF0ny+c4LPCT+HsvaSktx6NvTb1um984BhsvTtZQ7UNkybO2if4MnhrMdXFTky6axM0abqUo0
fXDqx/CsFoj7935VByvVW3jx4Ez4O4oEH1qzjzEiY3xowMxA3Y8/CKzi05AL29HoRd/fkbulYw5Q
Sy+gvY3N3sKvmBb9DTEqKChEZd6SkWo36e0WteYxy+VCtk2qpsCmwf2znja3TsbNO8SiuAVtapCQ
D7MesQE971Geyj5icq52TV5h5Xod6+COhlkkjqgGySwCVCrUMpG/1XM7IjTZlMDiZMlwDu0T5UJX
6AbiouJWJUUX01epWco+dD4t8VwK8bk5gcYHmv1puWtZG7OAYWGB+Q/zEFEsA5GEn4+APACbHI7x
XlUqEGGGuiMtbNb6fUwHa06HROHa5OZR/+52woNnxODRYUBCPgTZggig/0RkliI7aqOhL1RKTx+Q
GBrg9do83obeNCwLAGmujaUnoEUTEtJztXi42EPrjRzMESXbfhgZZK34QrJERAvoakOU2fis55LY
R4tNPoSDzspuwn+lq7rTleW9JB4l47rO6ntgpToFQr2uPVF1Zjbpp6AOQOQIk0w7Y6Xc6SS/38eB
/ntfrb2FOJjAJqM65o7U8htgBw89X9XPayrFrUsPKRTkhr1J9MPtuAGQnubL7u4xuvrntiGgRZwx
mR5iZ+RrsprCnHOenJiVcHqZzniKSmtgY+gD6Qn8wSKZgXQfRHqtQ13NQvybz7XgUfJE1CE/+lCm
K47XYcdSoJmfbnHRj0p2VNERGOBaTpYON49m5J6sKv1tLXYmf5/1gOzUUun8TGNci0b//P+DFhte
lZ2SVaxdhTvqN2fQjuaZaMEqyQnXnFJ4SLJiJqZuKtRoPM5FGHfV2Dwr3BeGGMXyUbvPp8jVFdK0
ageEuXONPlBZutJp7paQwrgxVxsBRXr3pYh761kkCwp5ITb+2q0vHKv3R5W2gIGaCkz1zW7Walh1
IfaBQhM2aoWX94nPprRT95qS14rlon8Ze/6GxHFYmiwAVbO+OCANiZMKdJgz2YVHDLtPJme6682z
uXuNqxTYIosT43zKM+NI3Nyt2KBxCzjroffI7yTi5MrVK2MMLjyege2DDaxYmOkExhPKfYx+B1JQ
T8CJscHxK+hGOVbSTLdNFxOn7wd0KLIdz9EnoM8u0tzbuuvipRtZM6P/Ex8GTxRyaxoDhHGFQceH
nn+S35NsnHGW86dJmQth+X2I+XuqtKpeJy8ShcBJgK2x7R2WS03rwOqto+nVICJQrlpPHIV5bXAY
YNbabhtekmMbR7xIy56mkwLH+fmY0SepkvpJ5S5ZfJfBBkiRxVDJwHKzfrwUoc5RzkMaQMW847Ci
N+t4k4q8XuLi3rZRoCz2GPdVDdc79ZPzmErbRAEdwjybSVB1WYg8nV/LwE37UBhgIjtOuOoRZFYb
+4UiqNpZ0fURaAo6ZotEypnvNEZeZFRqdjS12y65VBjxncjfv+OisJxbV7FL2LsroIRtj2ZZG+fg
f0Sg5Q7ecFH4fPiGTgexYamOjb3BvY37xfNHEsEi0+AeNHpRvv83hkiR6ffn4wfo8fkgLuyHZvj6
WIJjr5lYZ5yKMYcrvPtbm2K/LD/n1YHJy3BPjGTg/8+GPOUQUqzS/F+QOCzweWBiNLGE3bfnnmmS
60HGxrgzqDQQR6olcmvKxRwYTm22fupbmTEzo7MBdrzRLtYGZDhOFlQKIf5URpfqnGHFn1/c/z5d
1DCCTJiT/i6NLDGtAOmpjnlMcwDJpboT01Ulery1bBVdCUE9IUESj/ndlHaSlMsq2V76Bz+P+REU
F1OL//EXUUcaHx3g3FTCDrFY5a8r7O6GCw3CKJsYRYCItYzB7dgSd/1uO15chDqJyPzgSdVxAfnz
uxGg/c6WNpqvAo40BfGoCaHLMAT2Td5uCWYESYFVy/Oe2yw6Ek+u/U6l7N5JHZpxEo6ncxwr6iu1
1P9/tyHLo+gFTm9OfCDWHgv6pMBNCTxjzV4P+9ARf397mqVvnmGSB7RbDJ0Hno1OYLJKO5MyMlaJ
kfSkavvQSE4KcqgyltNkSM8PX9siyS3a5xv1OcZRPjJ4rW8pjyoUTWZxBL8rfAWSmjWzAXBSeu8T
MOKVFjs1lyHsYPUDzIj4Y/FHDio7z2pLgVRXBAwO5/pecpK18gRx5pllQu4opjc4k3mnCAHEFJPr
L9lVEFuSWGNs8nYP/v8GxOT0D/pPe2mKuD1y5qMA4ju6YahK2ugJdVzJTMarB1R3Spr/OTIL06Ql
SFLCAw2EI9AJW9bl56uGwvTp3qDkumC8aJBXtUOykDD9CXsqIVE0/XQSb9tx6ttTPwj+CaiSjHyk
FI8SZ75qD1AO/ylvfZiotz/EQ00y9gOSPotT9wy6+l3BEmlQUTEJTrQzorZa57zDj09JPZeA1Uww
AqKFqxGAAtJJ3WGIz0RATVzeKAz/yDe00VpQYlsRYIxS7pDQL16kodW9UwuO8wtcF4IhSqoGKPWR
/Jgz7BOiaIrz6ZvzBbPTwHI/rKMRBIBR71TZSBOhh7hJBedAkIxcIn567HyPHfsniq5mgcAZzqw6
SzKZG5x4U4B0f+pKQL/AqEfG0lLQuoII7KxQGYGvmGbW0nnwtPeOzRCI3yPu8otuABXHDOakzT2h
Mbk6dT7XjXiU/2NEBx2jrdAlEw20lQlX+ZzJ5b5ddBxdud1/98uVaag3Pg+gGxbJc/cUQS8x7Uj0
MfOcca64Poldf7wPFviUs5mWsPHB6gRX9U3EZZwXl4wicjPnsS6lztBu7SlOxUByLI4rNyfKWJsD
23PVzyStN68PrjTM81c6fG0PXCfen+DrNbeh4s9A0w4vGWhwgADN4DKhYZX0ViTEB/jy8gwrxZVN
DDOTddrfkeaOfTuIupebkzh3J2Nd5YI/Dwh8AqbX2NUiYj3LPJiBaj3s3on/WHbF0GgbixMjS0g2
gADQ/42RQjGvaErCgyo4YYZ+6gPs5obIbPCJLvV1z4GWc7zElnjikSJrPMWXhjWVisGU7QZ9Z/pQ
wRmKUmTwa5tH6nEg1ytzxWBaGexvYuqWXaFVPdIJz7UQg+Y3mf2JmGTBcalGqYBu1ZNFFyIv7Cez
xgXp4Y715xb8qWrHP18WxZ/xqubde9UJodYKwcYowl3f72cS2fj9dDQu8rYiqiGgq9rlBEqaXtJc
cJskfWiU6496Nh7C/Je6fjZUgMP7l3uyRPazKdMIXxSIumnAmDTnrwa6Udel3QbdsAfTEIUOr+mM
pn+uANB/ZepdC9sJjKnliWFOADO5aA7RK2/GUsvtDBD5x5/PTdfChNYH1VMUzK6eRdgq7fYbZNLg
PCQSOOOFBevKoCB/gInvrIoiKtHh06LXxgxPNEFvy0z0/OZwgDr/xxlUbIRqMSBzbmq1ZqA6evWt
7uPIIMxNE3gA7dGf1S1x3GHCRDY8oTtkJglORr9UYW4mpsGsL03/7Wip9oOm5hsxD+Idtlm0Cnnj
j5ymATCZdTmBSd4WlEwKN2T9Rrl9O9KPx2b+m3dwyLrs8/AhXVsT0l0yJsgfv9NadXaobaymvJf5
oAm27kLL5bCMNqAYesupDgo0dIOdbRynJGsVwIwRA1pvAitrHxC+W2ahOePtIW634lVLU7Ui2xXo
dzXBFcgcnKgoR3peQaV17YqxQdgkkpaLwumECtpw89PLTUBgFQXK6MKTq0za2Rf4UH4Q1S1dD8k3
3eJ15U0pPrk0iBNZ1/gDIPYicwuzmDfL+kYCq95jmN5Ujb4cdcHAWn3ibqRqhXAkbl722lf8LpfM
tOosDJmVQyCKJAkf3ue/d8QsLOtA3fCDVf95FfYCaQ1CYUp0MRpEBB4K5jQxV2LQ/94vlN93HclK
WY4P+paV0PW4byU7KyV12haQcbVgNVVIF3EQN/OkNKDZc+0+x7WCMRaCUWSVHD/c6YJq+Kipat1S
TiNlJjcsLts7R6jwLc0MeeF7L2hwOlogkUeefCaI9psMuQihixdBu6RHEBB/8SzMr940TO5WO0E9
sMhWcZsi79YPADMiEaLBF851qQzZ1CQuSpF5U15i6vEEI6Z4wLLaRMpW2Xf+eYEeXedilO6YtB9N
vJE01aqUcHvaDGX7oSIM3XmyqomQ7lB3+7mVkN+YbbPyjlNu3kMLDOuueaBvyWreHK6CSm1uQeP5
R3eXmBtNQaQraBSWrKwmVoX77+XMql+/01Av3uO27iItJ1fZabqpBfRnGpPSOO0HCoPHQe9K7aya
Bl0tRuYKAjO1pOyA65UlbmKq7y06cvI6o0BWGRgquv9Y8diFKkpERQVckfU4c0WHOfIw5FrS8Slu
mcEKmlxlAOQunB0lAw7jA+FPwIjhKeFQl8jQAdPWdvy+o/yFocu3byXcUSouWgXK9XBBMZphvsNa
zqPnQ+154I4+R8nyB9r/eUv47lEFE0FD41p96HCPkxGMBUnUulg/Da2IRXYXkFnRr/JYAIgYJ+IN
moFvwHbLZw/NtyVIR0H52YfDhlRPWfpkXOFfoHHfTmjdD/MXH+OPK1n/n6p5a8BiX3J0WR/jYSFQ
fubJHzPKbUI/zZG2p+JMuD3Nk2RrOw5RdlocyinufFDgpc7MM1PH+ujrpfPiM2PbU1Jv2eNf8G5y
cMng2oiYDraAj5OXP0u96KXPxnDCTpQGbVaAM6exYl1/jeCtv5P05mrYWniRaBKaddvSCre/13xH
+j/sE4eirzGbjIWMPUb19XFfMdEfwOpSBmKAvoemQisZzDXyDg1ab+mvofprQICwZXAnFJKKVQPH
BNQ7TwxOVq59fUeS3aLCxP/XJGoEqXt4m88WNvNGe3D97wCGI7dIbvAzZ2501Cu9PuMFtmVgVlOe
k+sh+1bfOkDdeyvKf6n4EY9Vfe7ikSRe1TSAgawNPYnVCyrFyoI7OCVCcFExrByhOE/iV5eTnao5
LJBDmygfCLyHt6mx7RSP3JR2F2OPmSM7G00AKeCdrkQguUK2mWk31c0nF9lPGah/Szi7OwE3OKtO
aAC6Pj0EAyS67hsFkUNzEP7nQ+cqkMzuH4HA4/ssRjXPv7gNUHkzRXq2wyg7vqsCo609Bk+XvizB
jUJhn7smDbPZ5rO0UPd4hd/6EKZ9UhHEZU50vaGWFpBLS+Wk7ZM4hdBrBcZ52TobhygUyg3QAlHF
jjn/tel3CXcq4LcOCw5Lyr8iLpUL3tfMJRhvDMF7BiDrZ+xZ4KeyRKFWBL44ULyWNElUvthAC5Rr
Lf1VRP68JcdOp60eZ2yTRQItjmWFB/dAR4+pyWntPXNwoJG3GQZS70N4aRJHQ0xqnEqMIdIaDp2v
/cuKUsFt/nXeubLqwwf4T1W067TcqAqZLurzzEy5Xzse/gEEB563zWJKzHE4Riimp2y+JL0VlGlv
F/XQLfT10/MrIrJBXW/4u7SubKJgoN+3aCuxzvOVYbWc8e5R2+TT/wzO8hO7tjOcBGDq9vv9ffxh
RGk7Z3qBL7qetcZanTyj6fOiwVfswiAmvTsvo1FxwXjQU6417oZouThtmYsW6uytOn/M0nI5FTpa
h5G39njAJ7o1gl/EzreH+a1u8OQG7ZwhiTHl68Z2xCQVUv1lryV0fI61Is7B8xh4W5s4Wxha++gn
XAmZ8VM4oxSurXxSHA+gmZZcUqwwVIhJlyAPmraCQnGrK2C+x1p9UQpiYsZfHlVsYIs+lhCczssZ
L3cXWzuOZi6k7V3SaN9U5umfbDIjrqG6Tfsf+RzoNQEpetm1OKMswKWufyucs5rtHmjeyx3oBKHX
Y8TbV4CAv5RZduHsnPE2UzlEkegp+9Rf5O+GZievh5Xk3bM2CkhzTOYGttGDGw6YQyCimtm7Fp12
/MgdW/nn+SJQ5DWorh5vbha/efbcFuvfKand+6RUQ2X6Gx2ZEwgKnOO+dTJuSGw4xepLFdTUmYcn
g0v1UPmOesvMPtHnLswOmZhSGeevwn3Sw7kDQ+za1e3k+yv7bdYsHv7izFHYrfay8QEuHFau7VKe
3GjCz0014KAgmIS53tHcTdlYu6u7swMSgUzFWvqdZgdgSntsCQy8I+T2GUGLB8Jk6j9p1F5byzME
X0KvkciFRzjXpv8AGpfgC0WSK2+gAHHpRAFL0MQKhg2NkIa0CEIZBA80zIAqNREhHFD+V0sx+9X8
zgUpkgvFqj1lKHL3gJ434F/maQt+6jyY6ZrC/IX1uPSMJ2riudSxSwNlGubLKOobVzVn4pY3yJ0V
ovp/miYLX0VpjzrGz81fiUQhXjuxD4FooCDSnxxeW4BctUfqAriQlm+D5av6XyJpdXRFNe1g2KG8
4y0Qe/qQJCyAnRTMw84UyUYSil2CzrrWXQA5qHup+4A7p4R7iRmJ5zW/ygCO1W6zrH0lhTk8x5CN
0gcL8aUNU9x0y5upmj3NuJP5WYGvhRztii6fKtYoV6Rhm13QXmWhTYMl6jRzZq9cBFYwyLm9+sEY
UY6FWcJU1/a2w0Du955G9KraGFbH2Dl8pyTB0q+EIvj9fXFIYG5r/mcsOS5DIrm5f3nJcgmm/7cS
yhfIJ7upQ5BJmqiDnfy6d8YhogPNsdiIAZ4CKotABZR9hmC4/JsNeX5rRo37nId9WQctuwUE5Whl
HYsC8ZRf3E1I6sAR5EEyH3Rccd7TeZRU4MBjCxiZe7LGqEEUaOIHl+ngyAleYqbfssRXVQtYdHS2
BIizC+9s2BfqBi1VSd4baow0SuY2nlOXdWneYmK+MHUG030ODxg5jDRLCAUktSLFPH2EWHkSUYNp
g6YvfCMWtpPdm2jKNOx3ofKRhib+0ffhzs0PYVbLK0WIzMume3Ou27aTD3VqSwZeaGjIG7gNSehE
WjDlqN2I9UjT2D4iZzyGyBMKnuOGC0ddbKDX7ww4DSsoYnoGUlvkpMttm5ytK2o+iEzRRVndgd19
OLWiep8SlhtBhjTbhFkxwnATeJfBVI8+zpkQY9SCqTC55rDeWHhP0n/32CP1FkoNFd/knTrJSM88
rHNg9ZN5r8/TxJ3xb0RnMKhTctFyLT3ew4xtMrHNZHeZLXzhWuuwO8IUV6RZXsj3VSS0MOjZnIk1
9WmwIe7ioWEy66OfcUw+9mf6THogbnSxj4h6gWKO1bay26BV9+x7HKMgIuDRCG6B6uqH1MSflcsy
SpefhlXRJZZlZQGz95EV3vT7Zyl7u88MREO8pQKTJ0Qdomnf7ut03L47pSHvMgqrKBv1AmV73Ejz
l2IR7GyxvkaMIy4Wex939rkb0n/hcyWRdGZzrcTY7rZI2e3ldfQuuMglcKQAf9jtzgGwKDq44TKZ
e2ndk2QEo8lr5nwNNbE38AP8x1jqEtqmlS6d4MMRYfkPc4c6fM8yOYy1QgFWPPbEYW58AxVpBBK/
SCcW1FD9XF38IWnx8KlT0mSFh7OM3KcHMCmJJb3LmmXe9jLCoQfdhw/dxpvv9I9TF0BIU0ksF2MS
wgnGlYfD1g6JV3AnB9amph2hkExCk1CZsURE8rrYVzuxT3LB1QskkRhCXOdb5lRfo2+gnDkb0DoG
rTS7UytMRxP0exQmW61td1uDnwSLU3spJaZY4+NmJDabf9vP0SXeSF6AGOLPROAQ7sLbpqawoejA
X4Ja4Otko2wfSegCmMKGcucNgH30bqx6RrHOJGxuRdWB/iqx3HWGpszBWCbD0G5AFX0tnJLOGChq
5M66priFp2d2kajWsALcw655Ev4X5QNFT436MkHmDX9TzRZz1rNE8wrg54K7buNjVcFw46JID1Rv
qXw+aOcNuNK/TMQEEXCDZh+osTP72qrNkNLOOZEXwEytCDrEswsxDkgV+wF5GcJGr1pGr+o6ufxO
cDuEWHcPj4tNLuBjMcnX9PI5JzdRPQckfREfhdtBzNjI3JSBTEHZaM9iqGefCAJKk1E0bAqQ3yxs
xPMWIBDtASNpFoFDUYKff2iiyt7MwAr2Z5Pi/uZJXVkqWJtt0HspEoiZpRSYpPWTpLI1wPyD6RJh
b1RrfOEadnj9EJ5seuVoxSW/L/4oZa14MBzMFRQPOx99yA5NjNQcb8Fncpgx6UvtpvdicEheYprd
qnx1ZpfmeaXth3q1ftk9s2/EcOxT7mjoYbFuCPXgBmPSOzr7+geUTkMsMDIgmTWntEmv/OmzOgrq
Lxv1O1wdceEuuY60SUCUrtv5y2jbk//m9O9W+tMjbS06awSGwpNWk4QMCiMLKhKWEkQYTmQM0bJG
SlLJlyhBxv6ymrFWFeQ+iuZ5Q7xu0Gbn36KT50Aq9gq4JGJmK0fjffZiEJh6looMpEHDFjGRpJuP
t1TP3pP/gHDzweQ/8V8ubzt8CFxjMDHwGD46X+MfGemBJD6ynnNv2bxEwl0JvrUS2DlWdHt20Xk1
h6QJuvdRIy9H10GEnpIOP/ZoI/kocpqCm9NcfCFSbsGMXSL+A6pHykI0xi/3asJ2MoQvUt1xvqeT
vmbz/HQypOj46zSmd10S4WPRX3R4cX94EmcbJ8whNU/6gJujJppD4hbM2Jbk7gizxd8EgzVKuWFe
EP2Mf2JysKJW6Tv134Ft/vRJKXoH6U+xKQLupmnKSYPTtpi+Zd1qEoZb6BEq8F3HuAsL5AG1HiTa
dx0/21hIIz3pk91xJCWQYLSTujmVWGvglUGy0DSKI+WRwFzTTYp/arjD52r/dvrkMNsB+eXB0GN+
bsMPutwO1B0CWa1Z77oaGkHMe/nnUhpvq2BNMBXx8ZH8Tx5OdrmcyBu2A0EYzLrx36CrkuVmnVUM
iBqN0V0FJijk0r70kgmH8mSrPE+q4aU8Yogp5uHqxz7taaSSZ74MJKpXanbb/jDoJ69iraE44prr
kydIKOqnaYLsRTjiEy8F7Ws0Ib4ZNrnOc6CWAuXSBbhWJsYFOUqjUCxsel2GQBvrEDVvgl6ve1DS
txg45YqCSHxzbmHMNhU0SxEH8Em46qjBHOCre5EThx4sF8lXSbjah+Ortnr6k7MS0tbNn2Oo8shB
1NK4fZkGxxerBiIe+GD7DmdIJ++N5PP/OOhcoJEDEFZdQxnmnSEqpQWOe3wo2jAv8cTchdg/3Qzg
qYTVA4orxLo2+c1rS642cH72QC+0yZePKjxYhfMWGQlYPuxkFEqOmwWU6WJw5CA9JbOxWomkrcVi
fewEipQO5izsTatfx58hVV56R+WE2cI+HNMM2QVxHJmYBNvzyN6Cza3aEvfrAgwwB2tYFZV/koOR
QHZZzbiqpiQzjmQNscB5+2ISW8I5ZJa8qolLBHAm4qyr+NSfBin5170QoyecAEOCZy15iVIX/6+K
G3N91pWEgM5YaKpA8OFCl+Btc328WjKxnw+Q1p1iYPGNQ3HCI49ZrPruWm/gub6muEq0Q0kUiHzv
NWGIjqhEH4zAto3H53FvnEkuKcD+DrYUyw3iYOTI3XiAIdANMu5Rpft+WzpJVH/KFHVnck5z4FOY
nmVP6vZpFU0GLjK9T3NiTe3uDHBUE3GEy+LM4NdfBTSFizMkvLQ+ujiGGbeWhy6cpB2C5bOXNVbx
GCSo+c3xlrbEjgpnkPnf7fJ9JZsp5jfDSpaPCJzUfk8QxXEuIwPoHxFxfJHLpdE/5ntxzCC79BOd
HWWE6qTN9B6swf2RQyhwjnDHpYkyZ/d3WtRyohIleCKuq7gjQuoQ0hpAhBnlQi6GE26Aya2/9b+T
XfdOMf2QnfGAhniLUShiQWOhMlC41wkoFGT9kV59CFxmwnmPJb6eplbH9LoBAidAqr4ppLdIBgWz
UokKls9gQvSGrWXcga/TPyBZkg/Q/VSsxg51OKfr/Znf2cYy++AVPylp+7gl57PKfCBlnqW7Mpae
3cfUsMBkfdH7UZ3/5JE+MEUK3DLIk/r6Zfci12HNnlwn/guQA5Y3WbvAgvHXvPSiYtjDIvCwCShI
ODbksPimw5aY7lUH9DJp2aell8dd8rWqSU3xjGc+/qtuTdnjp9DFK8h3UCQZyHongLc5LeQWS6Fd
lN8GY6YrNivaYOzHkW+TbXL1O1WhkhJ/xxG/AeCJgBvtgOf3QQS92qX3Ucqz6MbCKREUS6zPmmLw
205B1ZAdDZc99dj5iguONVsvj0OIEUDAwMLZ5PLfIGH9T3x6XDLcgx2I3LB0UtSx1gGDZ9Xm8sbk
WYSdVXCor5omX+LMcEVzZqduMsn9N/cKHHmRxYr+Ul7/0zBGYakhho4+o5k85ZPg3/v5L4RUfUdk
jWU6Ev1QfpanL5azI/hAzPR1Qfr7zz4pgRVaKr5kMUy64ySh3kGM5GrZDRFq3kujzS21CrNjBZHe
bMSAhMq1H/DBHTSwqVTWRhHG60aVB/TzgndBl6n7Yeddlop6v3RieDRioSHOALGNDsksds4dly81
e1elSJe9FkxeHjlJouEOQpT4KilQ5Oq4YYCGGiTXdZsLJ/lo+oYod9kjoYi7VuDq5vSXjUgU6DZB
Np0Tbme76RBKn71oK2kPJ2PXW0UhpB7YblAZtE6KFS86GIh2Y8Vm3wiV2+vcHU1Wn6HHoiEloL07
UcrcWunZJ7ztVSr93W0tkZq/tapwLnaE+TLVp2Piq+hEOOD2jayMk2pmBzMK1XnR/RWIHjUpPTFp
7wewuuBg4B54bPp9BEA8PU51LU6kmjTzoWyYKqdXQUJJSXq0wc1782Sbg/QwcTtEt/asK/is0AjH
7gg9OPis3A+gjthHVFsv0nnIHdET3rfsriFJsPoYY6scJGz8yHy1sRrx9M4Td12TTiaKXJ63zYB6
q9JEPe3jDCJjI0hG9wGi6p2jOk7d1AIY7vsKRLpNolzffNEbv0emM1VkGJyIWOZ0Q/uqydVUQu9Y
K3nU96oU1vb4j0FDAXhV2SlTGdhn03TEfzAc7nVZZ7WNFQUUm9dlcuYE26mIVumoGoOqpkWGv2KO
qNV9cTf3yJkeLDu1BlwbpragX6wT0Fy822xZ+haS8T/6CYo27SWLBx9dv1qGSqTTfK0h4IUIUFJW
1rkG5ducp/CNcQgDQjdIVQeZ47NxkY7FNEeHdIbZrSZ3xA2A5cHscUgXE5vIATwgc1sPRSRGnKhI
0MoZ9s0qkOM9F9bQ+cRCnRc62FVi21ZEKur7j/TPuY/cnhxTvEyFmAnaUr78O7Pn7Ml8FIGewl6J
36750N+HnpPkMnGOwpx3UwBvmjL+jJeEAVVvtUCTCpkYuOdF+ljEifa8gVj/mNarRST2J7kRVXzR
gX7829DCglcwKX4Xl8KI28z+MFke8GN9BKmSq09vJ85Tb5EVMz3zIuEwhIhUJ4wiJpm7fBX4Q15l
jmMwXlAeaeHwTDmWT3wa5dbImxiRqa4b70YrvO6Bx5bwkJ+5FSPXgCQZyAnN9Ucww3K+vmWi6MO9
J/QJssZ5xe3jDavqjvdV9pxqZhzSlrDlboaItxXbcbko7zLE29JVeBj+/fqBFMqMu/yLtRiy0yBh
7ng13LzEMBOlt2JmpnOpJhzBw4ysSSDE2bGwVNm4RkxkWDnrrviNRbsfdC87El7tMOnIm6Fb7Uty
kELEXzSi3KhUaJ+jhJ9aqH0uXiodfn/iy289mlfYwx0gb4lPmuYzXuca/+kFVO1L6Adf6ROfHNNl
sW3BLV7qEdo4h5AWpkwxqE5AeDSMQWWN4chZy/znjmrXIm9sCEF8st7FNEpleWYJ5bCJmpNQFJaQ
kRilwYB4rgvmk5N25Lvx/BjKOiGc3sQWyEM+vbqGN2ne9BusLltai+c7QVzhuRf+OHUzGmWZdQVs
PdbtMpbXVW25/xJ6CuCfPysc+wCM5VtR1uS2+HQimJ/zyQKKROyZUnC8nNuhU1P3ifjdJ8Eoe6H2
qjIpreKr+Ax2Hb1jgBIX6Lm9ldemaVPMrSbgZYGpmxgeLcRIKmsjtBO7PztwfMectj8tbVeeJ6UG
+9VL2OiMlxMMNnxZLCTb8XPT4RkCP9M5qW/C7TujMZ1kZELTAoI8RNvhBBYbTjT7jjkj+hIgSjP5
/TwyN6ehLKCom+rfHpGonZQTy32PVsWuUbuA0kdzfiDwFO2TbHcqqv4NHXE3CPhfNd0U4/XAMj3s
yDIexAZvWBO22g/CxtpxwKahDmQEmtIwBq2BAfyXYm/G0ljlKRAuxM60W9xh4z63mNMnWLk54rG5
Cg3XfqYCiEmTTmDUoKv/BCF/9XN4uk6SIVo5+WSUATjVFUaGjyWasjip/8w5P66s1AirA4+qu8yL
UiP/15ys9vU3RNz6iIbX9KN7qkQdP8FL1hn5p8VdH5BNKkkCoe/lx8D6FZ3biyQrePHRwa0iueXE
LDwGWr6igWBW+kLkuW+oOTaqThhSeQoP5/w18DwhqeQf0SuaPsFF2cUQ52WwPmNLzqLb7tygx00v
kG79Xy6sypln2Da9f8a+c8Xud/hwCtKPX31gVjc7V5Dj7bbj6Z3YZ4fmKJ6RADiLWni8xVHgMWwF
zqb2gsRxqPBEXLj1vwFJnhJwnaJow5LsYj1GmXZ7uZKx97lK6DJ/IXA+cU0oVEanlSOrN3zPtq9m
o+ZoWZWSM+YMgx8CHlfIMPakBRmQffVPfga9uJHZx3dWssJoMmC/Pwkl/FXbGJf88mxkxLcHAgLi
L+oyh0mYwHmH3D/+NDwxF6UeSOkHu1JPrrulQmsMzQVHAMnEiXF4WA+vqyKnd3xaw5EXOILTN76o
JLxgEM/4eO7Fe8X/U1pzNBtAIZ/iBq5y3n9PgbUprghnN5HfXhMjeKtPOlYnrF1d39+F7iyP27iJ
E4Tl1d0S62zIPqhor2dQfFMkVcg5u2RVgiQmjAc5uervRp7/BfkXkBPwmZ6wMxmWHDUp/xbzqlMc
sYOFAVYpEkObbfKapGGvYdqhbXhmDaHzZ62GyfhWFBEWePV7Ph3h0zF+9qIb5i2ZMgv0zjBm+D9u
nEJodm53+JNw/qmlQwvKvcvD7KK4skSeU/z3+xFwS9Vs/wcSvtdeEK7NI/w5JscYn80/w60MPTvM
tSohkvHz8VlgPoBLS5NOeRe1e70YUfZP1MQrveU+XtkZ6dUnGEJAtg176MmNjtG7gEJREZP3fsLN
bqX17HIeQ0M+MLkkIvOrtUtHXht9qKOenqFOkNXsheCIzWfFpzRN379LpiiivYoOKCTdlXzHB/c9
0ricQSh8UJZegfEQtldM53e+yqxLDDy7jUEYmxPig4H3WXm5bw1g0RUItFmZEB6enkcLYW+xqANC
7sJrbygM8RESj/InFWj4aWfSpyis9aXVwm+t+9AnsivddRTg6Y2cgjbN5D/vSTqa2vloTb/c4pKg
m328JOoAq0xNTkXnIhBKi+PXEviwKdJ+/1xTkg/kLDttMNx6xW9jtli04ROnDVQzIHK2r/GUXkjq
kRtDG8Yqc/SVVlwWSl7mxVkAwtikHXCDzPnCtyL5mPtUV3Z9NXl4KtNMofkBKszAebBDx7wh+DkO
UCEiHIunLMtS6vO5lzBvzglZ6/T+LvmOYQ9OXBLZPPt3j2MJRDp7xliW3IdlNAi9lbFhxM1o43T8
6BwxTwefuUVJJBwW3wHOrmag2XiLvg5FKZYKiNYVujJu6xhHYJejzoXSZkNT/szrUnu+D0W3OOhu
xuLPaIh6il5/SGk8L2jW1CQGnUgLDUoaJ/FnzdrsL9m10F/JaT2uVd4yD6g5bomPsPQrUw4J6VID
cXyOC5hP4xNswDo09Ymwi7OkBBPHz9V9UMjeQdxSfNmCziwWEEDHp+MAbTEu9NUp3sQxoBtyMeis
MULIdopTNUm1q4uKDOefVPsJg1OhOi7swCh/5bj1dku6buUNjhfiz/m/RBiOpv0R1b1RYuWzBe0t
b52mRhXoUKqF9+pJVKDX1SGIf0J8vmJ/TsnjycJyb1nSuqbbMq+7oYsmcYs4c8HZLVUMQlhjCJ2s
ZgWygz6SnXnjYjlzOWzek6tCnpCOdNVL793ZliFefDXgX2AxmqDv8g/hn8kDdrudcqwQ6Qgutie/
jgVnDGJ5H0L77S7U7nYsa1sXrDodhfcQWOvTGI3y4/neG1Clsgrfa1I24FoGUvTkHdUUOZtiahiw
6uy3x6ujU38Is9Gw3N3ZIHkzgaKmhtl7SYCS/5Zz2QLgSLhhJ0t1drOau8ua8MbLGEvRFJlggVFx
/Q+wj7jI57CwXrdI4gfa6x1kOKpQIcQmnYl4oHJSqT7Y6PdUAZSXYXJwFwM1F15MAlORUCzUQFeh
i11lWN6H4PhnxNeS98jSmRQpMRfQdE1KSb1WqwAkcO8jQ5DFW+blLaGNbXxUTGo+YL0tAwPq0ZHW
HE77Tyl2tJvQDQGar26/1j1zoB/zXPaJ9WCy9OGTCU0Jn+XrMeHBvRkUXnPKLkZSWWRamixOBjKv
IiyoW86VggpLJMO1eabJz6X0rMkCy06Q/lhRvcBnaIzkUCgx1uSS4E7HFbEyk6zQawO38/l5kW4G
2k5dUGYPPvqDsQZ2AXnQoeeTHfbNHvZ0R/NqbHT/k1xiK9AFtt8aHY/vZ11g/96y2unjJPD2LseT
dsljGOF0xHlbtHW0owFTuZT96LmQxDOR4V1D6057/ZTxqWzzOS3KIWEr+TyMExKxCB5lixHdN1vT
tvkfSGcqVqkrHJ8xY/JCyBVtb+6MmW+vTirqAFlNhf2DcRTSUL0scExQX7QJPkvuWew2+feaoGF2
5HGLDv6YTTAZ7DlCh5ndczRlmuK6YzWoQjfao5SiCXFcsGg/JgFPpu1XnlTcULZvz9t7UknM2xYQ
Ua6ngFTQm2VCP7TRfL5cqv4P/QK1KWtHgYRtzDVja9cjxMqhQQ8mtTTiKXIFRSvInTKzkQYgn57n
kzl+ySHgWgWT91CL4uURyPi8bf9IbF5M31X+ddF6Te6ZQaleX2jafE7LQz4e+5D0wuhRGaVamHcR
w31qSSKq1IaXwJiezmr3pl7vRJQp3+kLpPYIm66cGDf257xHgiD3sbRaZ9tmiAVkXke642lvNAbw
PmviIUOCKswZGCZMFkAgDT4Q35b8THhrSliYsszoJw173LOjnjAdovenI4NoWW1PZSV7TMDfDD49
BZmduzHGVMC/Zm23iFh+q/kfr5/GTp+gw8i7MY4QpyY2KcsrANaFBgTqPit4GLH1UFvSSuB+JN12
DN89UhyWO2ZcVTUojE9igZBXL56ClE/k2vrmYWQ1NXujxaSAD9uyrmiM4AZ4HB7pvku4PLjCGasK
V8NU5muz3VnJWkXFtGH+UwHhQTTQJO1uKLln87yONhB61tYNev3bYtcKkqgl3jc9V9d3DndTPK9B
iNNlpFFDtxShdzVufTG8LDeZTYH+GP89fnH6PA0Qei18lq6up8FrgWGd6K3N7BjZcgQAC60N43CF
sUswX2vYHPqteT1mgU8Gux/48ogggRChVIa/R/Dy8JWOASVwKF/Wj+BKJg2RoIlFpMIqxInXUVuQ
DElesKd9bKa9sC/6pqmT856DqDbmD5R8CEiTGBqf191C2Ztj6M51ymOz0cwyOS8t+2I77NPmmf7A
Aeom+pnVXjsJ1ElKz+/RbaSEuXanaBA387/5l7yk9MrAAP7wEReAfEEO7mHRDeMQ7wfvHBofV5Xh
2sZhs5zhlpMI6fc7GATkNFVVPtaLVlhwIZEbsmmjKW8I51Vzl/u/fBpzbrer4PZe1li3PbazQTGm
rEm1lO4R7qUoAVUsLhElv3AdS5SV98T9KbOBgnkCF2o3njt4GtmDRFY9rtcObJvXbL8svt02adPJ
ptXHlDuAl0Mts36g3K9CY9LoXu43nX82IDIM5nwq2lmHYAp5DFEUbtreArwKS3gnhn1vxR7HPV04
Q9VnjO6O8fp/00xIpqF4GvzkOMeTM1B6gTDG00KvdI1VXroBLF3QxJme6J2sXJ8KlcDR6nacVUyq
4VZ0AWA1EX56CBRKXL/fFKX4M+eTyW4BTc5dT0UD76U8cGpAsYHAxaRhW1Zkf2W6OicgWRk4yA4h
1eVEdjl+dcF87T+6vfqaLs/0rvlyh9JFsPsOMk+4LXee1mMxOrS7LPQ17bSzA7BULvMDqyf2gHCR
1i/Gp1el11Tfcqf6Q5g6isVLUStoxV1uMUMGRIxBxvOhRAcohunKZTUQwPmJPHUZnWgmZtyhyheA
KCR7UxH9zHZ/ktNMeqHQMtDTfGDirL+zJj7oHvZ/mdAUsdtahZYOW6otXOdVzGHU9ad6FpUxoK9F
a7xfM3KZhYhTwMrtAeV1aZFyarY9OK3JsPNzRVSVFf5OFBd7mn7FlhIyEGyyUBZUznJPh/doqkj1
8vqS4E+yHRRPHy8lFl1DxWp9TKiRAEzhGYK+PTC77EW7uUzuGxwiISRwdcZr6nfVbwiM1a0GyvNW
fmU020LsZoy7DVCSGNGrec+fwkrQhkBYQxP5PU5dhyr4Qu9S2VJBo0Ikpr+GUZNQ/wrFnCXofBqZ
U4a7vrkEFWNxUnys9l8hv3QNTrqo6z1mdVafXNkEQ6MmgDuVQ+41kTRzhpXdMvrPnxS3zOqB/ZHA
n2UQxgrk6hphBrDy/3fnvKcR1oqjurfyWF/TIEHQHggIzKtjhV8tiVC9EKjyamDL9Iex3BFGipnE
xAOhYOeWgIsTe3169C2e007leFBByZhfCV5s6vXdx1BVD3Vb3uLnsF1eOd8+UxxKASkiVV/k67+r
YBfUtU9j0Iq+8YqLsgMi59w1bs+3abIg4aYYqXF8ipkBLyGjgVZJH9DO+cuFSEdcKJ0MnV2C3vCY
l7HOeZf/bBtC5GCkPwZtvB3mEnKNFyIkhkZ+raNN5zU9TTnmdDuRveNsv2KOY0xQ+wIbwtxxSTA2
K6hJxB+Ou4W2InaEIE6wLqQCkhEXKpnoE8AydJpiqDmVcgDiee6zAcaxqy2dhnIXgAAdpuaL8mGZ
PbUpq3VBs1NH+aqH2kdnUa9lv6YIJjmnirRdtl0MIaixorjV5q46y3W5n2Ir4oLHJL66hPCxDDzT
dpIeXV2EG1xpNm8/KQ90DRDiTlpzy9Fe/mBAZ7EWp6yW1ME9SPej+Q2SQpv4YX/jF4Hjk/gWhs5g
JaSjNaZZBo9p27SNuRTf77nM8H0+wozTvS5U3Dg0o05TZjER1cgMiiPqh6ExJmc4DNRwztjuEDaN
k6aeToo6iBSvhaWI7BgJRxGhwDrkOXtOYjoNjdhQhDsyVA7sf8yb6uCJrlfd9AWX6USyTeYC132G
lbhog9PFc8EXb04r0aGYrGVyolcQyjMZMkQzdwMtzEGeh0ReW9djrsIP4OaQwsuUHivCDdMR8hEp
O0MlMbZTgh0cfMU/ratQePAZslebq1iEzEP6wP06O+1lc1HC4rG68f/H7kdT1T/W5JtwVHACHjc9
zuXOxUvsuSAl1sV9dXJtYnLzUj91T0ZZ+P8i/mqI+I7EeXrYE7NNzJrwRI6HkvuWJqgB+K3cP49B
+Jw8IECNtl42qWBSHX6bVG0CuEK5oZ2wQFyfrHvPhAs86lmwaYutSGtO6mkrrXLdsP1eSP3WtqK1
FLmlqt8+yW4t+6ux/wgmZfAvkzbx7zbViAzFyjq2OWyCBrkHNdnsIrWz1C9O4+CR/lBfuq7/Nnw6
rtJs0FTrcF9a0R6INS+Le10+N2N8W/jPcETwW0Xsiu9oqD9K6d4sOF2+YDGeXuWpWIJs2X1GST4x
iWx809hPzHxI5xtD2hiF2NTdj5QHOhhmbpcyt1RC7tqs76v2d4PufCtKruG2975MZNSR0GQhUREd
bH1cZYAGZdhZQAz/+B9jzC7piMD7jKXn0NzfPu88e0BsBreOhOB5++DRnzEROREZ/sFISSPotIDS
JAWVkyt1an499ybcyJbA41RVBikG4oCni7hS5w/4xWxhVxX4wr/M2y6iMhek+EKWqwoRz/yIFdvC
bD+cSl+y8UOg7XHBJESv1FwCEwT71qTfETTIeZ7r8VkGw7Jk/NATvbDaPEn2LjwZug1X+6w9y71a
cAc0tVYgoRKXIQG+x8OY/dPz5OwBcYwWOXh5lYnlpTFtbIG7n8OOYWRqunx6K345Ltok+Jxkoq0W
3AOP1oovQDGbFh/Z6GDJtm0wNnMwXMRlsGMn3yVsi2eZ+WO5vXGHhC+kDn/HgK2W3Phm9HmHNC9z
rK2PtJQIfUiUtDR29hO1xi+8PaoyOTrZaerS1+bwZu0ygtJiykFEkGn/vLrXzbVNWwt61SATsyJr
+4uMj7RHSbyTwqbXtvlJUuGnPJztMhhLiJVMKFDfcDULLp2ii7RelB7F9kY+gIHDJYFk/IGxr4ol
x8+F0+SiW0E9DPXa4tGuTMV7SaHmOjT0eMyK1GWgYBx3RmYD30fup6v1IQLzMphTZArv6J/jTbFq
6iTVuyBIi+4blb482SN3MUAMd2Q76FAS94LB/XGdKMdeKnxEQGHbTzVJLMFI1xZxirO2DUCpS4wS
TifhYRY8CARGKvQi5fsNXXfY4jtUrFZCqPvVt3k+CtMAV4WoUWWCfxYvL60T7mCfft2l8J4f9qMy
fCCY0eUDAyZkcDkkSXdkjfXGhOE+ZjRC4WorMGenYzeHbDqCY3L9L2Obenxqr/QbZkyCj2U9LgnP
PhVVO8WLtAmSLL7JJknkovUQxJLbPe0udUbFqne1J/Ko89anAPvTQIbIYLP1B3iYpXYJAxrSK06D
EThHv2us7XNtCBl/NKf+8rhhpDz2moQAI941/PdyNhBp50LF9M3zo71+urMWz6A2eUenDVDKQdjH
qu9crnH71ZRHwwlgxj74wGqxNTjkes3KsaIj6DjgesTuCuZhpsTBPqNureeO0oQNLBbWeOGXd75q
cpg+oqEHxOojPHkb6bXZPR8eNMxB++zV4n1PPpeY4JtiMhBSI2Za64skF/1ZX8yOkmpjYPTAefOK
kuaUnT7AemKnoFEf//BpIQvT6XjF6GXHnQJ51q43uPpNg61ZQdkm+wm83uJU1WyEg6Ps6tBGKZ8p
YjYDglrVnNf85uWN4GBPXgxjjrjaIYOvpjY8MkgDHOC7C1Vk1RdIZ3YmKkxqSnoS7cFfSX9PXxwy
5mSMpz6puI8dRFjl1V/HxvbNoIRRAYxHZ03SR2XRUgV34kkGcVLcL0ZZCwEvikQ4Bst1TDz6WV5B
81aPHsIXypD7dQbH+ZeelRMy1W5RKLeY43d25Nro2GityRhJ7a+61jxFwJ1SCtZXr/P03XlqvjcX
AbKujOesHAGMkYCk+d9q9HbayzCNMwyzSpjaIENU4IJPtM+h+BltkJZunbwvI1VkAG3Z0B9OhrzH
tUTStLuQD7PKItdBh6DKMEa3uyI/SlUuAXlvIpnE1flFaKJJL7Nl2sn+k8eOhm5tXDmVMmjDKYok
2pH3CXKXUhmOTFhoLKE7xWWyrBLrF7RXb2daliA9837dCaRuDUpSdR8Dr7nd6eQxAEbU2lZTLVXp
ud+diS94i1B4byx1FoLzM7zx1V+5aqEOHzXuLt1plslOYnvOJZOHOx8f9EeTCXI8TRnkXMTpxcSk
0zFBD5NUrKgQJSDya5nxmmks/flSEHdXQba5hWbLqLjxScmeA2FNQtO+yicV7IB500+QKnpT2ty5
i+9FQdsWF+LJr89pVLUEWx+GjfriRYiYcpLLGgCHaqYCmn4wZRtM7pa8k16hm3NW8xBysv+jXpQa
ZAcnWExIGXnwK2x25YZz51aFn0wfGYhy/kVI5eyE1i78vUE+SXHllPSAocAhQ0UzX1wruZBmO1BU
PmPB23wR1ISpOmlFdRfMo9UDuKTxLJMXAa1D3eIexXlUYFo9KFYZ+fwz22CLkUNfJTBXhtGWtRys
9YIho2zQ+/KwjcBZcvCGZcVW3lkzRZVsbR/HZiHEpstGIbQTwwZQyR8VTGm3MHNPvc3v2gP9nYRQ
D/lsJDbqxNCC19DsZN/w9SzYAR9Od4jj29nG/tBK320dYizQgBabiRD/I4xadhKWPfB0Y5XYwB0B
4+JkgTncp4ZXsGrRQJK8Ms9Kg5PIyimPb6EjdPVrl76YITW6NrC7AwwMB9dmatkr7sfPoeE8uvsp
9FU4lyRea02WUwn9w+8K7Xp7cS5ofiGG+hBa/PdMRZCRqDU46WJkszYxY+hmLm1FAsFrQ6ubgD3y
/Hre9OBCrEYUjb8fpnz8w0Ch9ZWfMYdAUYcpdtF4zB4skPs7P+hJOvbQHLGSroE7Dx+spM/N7nkI
wi+V7nPDpsbPsCritJkc6Fd8isvjG5q7oyFeISctGISrYlZndmZbH1QaDz06/UtFgDZ69t0+XMaO
8yLczbx/k9qEKOI7KKfHFmBhpkHJo04Gvtq9gBPHyD9XbeqyG5bzttg/tdkBKZcVFK0y0R7zxe/1
gjT02a0934ILuaLHpFT8ROp/oWYsneDXriC/U2j7PcxStfRw5XNoz5j0/fIji1YammeWgXjMMErt
ptOT4qDOpYvjJJrq5fOgtHjqum+kXykb8SCKphmdxLddx+Igqxb5LXm1Zyx/CzaXqlE5lQ8hR2vp
TpGchSVZjKFLdMTjj98jgaKdNMGxEDjfuWriVXC2GpxYgtmumOnMmbxf0mW47Qrl/g3Vd6MfIOl1
zULbiH4nP2PGASdyPu1+7uI3acd6Z0ud//fFrOQ9NpF/FKBM4gkPZpwga6y4d1quYriz3aD6H3Ie
b0ju6i6339GjI6Mz+ZnLY3jO4krcC14D/JtJkWHqe0N6DAJHtn1iLK07lUouJZU8zGfSiYoHbPI5
Ulwd2XV23zowOg+B71y7RqoZy+c5XsCv5sKYcUf2j+TbZuWB5EhucIAj6Wo+IVERSIOnBbaGqOlO
QuvsXk3hW41R4CnTofEEEDUXUjU8eAfLRXJaC1S3VlL8/BEEpRDxnAte8S5tF+wygpdbCe4Uoc/P
4+akPbkfW+FM/a/FPQ4nvwdrs3BQ0mt0jOwGSKba3MoTmBBeDXmyB9TrK4X31cC5cifx+1hxDDmW
wc6rqj/wbo8/piqSWB/feQ0A50FEl3C+MeRJkVltPPQdqYtFJHTh0FGy8dtk4rQ4GvcR3rncirY+
bm+dtDPKp4JHoECuA2YDVKGpkmH1adaU1x17y03PqIFPSszASt18NvWPrzRYpVGG9y7bxpw441P0
3uWo/0Sq7RBUo+SXIEXJE2OR4pt5fCYsQ08+iWfy9nNqZ+2jxoyarBKk5wCOuIpFll7uiIpHvaZi
mXmraZWpNNq9EuZBxYYHVTq/l+sSEUIhLX/RyCMEmWEV5dl4IEM4lbAkq8S1XSc5HRD+cU+7LiL4
iJPk83eQCc1/wntLSnIxV4wYowCB4q9rDY3OWet82w/cjjgyrKlx33O3M+F1/vj/InZm1fEofH8Q
FCl8ru+EBWr2eVrxNkTV6xVcv6CR5j96biAnecqXXsxxphxHLVgrt5Pu83ueYCQhr9qaykn+Q0DD
DyHjTYokajjBQP+LlN2AnrvaePp074EKCTqLfz8piB16ZSLWXyKx8eM5xur6ZpihpLAlSoH9lEJA
RlqMcZVXff+v208C6WQOeVIaTnVJ8MZR5cprx/PVeNEKDqKFlKR1JXoQiayFR69HZsl/z2IhseJt
iiUz8ViF8ohwhDnmWODOAfz+n87hNw0Gk6UB8lvnPSNrGCo3Ud7b8Vr6eJZi7Th1G423HX+Hhq6W
0QEM4CTQgVYO3D0m4fbLIccQ1Ndw53nYfDAcOQcYDwkob3x/XuwbveUTYei6kiLirQzqJJTtpjEv
RKRxR404ChM6Nkw5eu4tOT/u3dudSaZ90wkA0ohmkDTXdF4S+KG02DyR6k92YSt2KI0tXnzqCR8N
aHgWCp62MGlVkTanaa+IlwYihva3bZOgkcAgrf96QiMFv9h+381aMCkR/nfle1dtNj8oGJaZdYFH
6VXcfgTehNRVVfbY70itgGxKt1E4BN+J1J71XrYYR4bjBfWEVr5blFAG6JKUN2bzrdmu3QZrmH8w
+Ts1QIFp11w5XNuShXl9cNaQVpOYR1kbG36KywdBxumCVAa7G0A602UyZoNN6ypv6sJ3rWbYpiEV
lRhBPpp8TM2Rz8Ld1DOom8A5LSLsXrnVjPrauTOWPQY/jMW15CPHTDPj21k66tZKbhlUJEgIb9dz
O2wFosRVtdX0otQCE7yhj3iwtXJgI+ucIBDZskkIqK22Gx4EmsAREEZuuBqw2+4WAji51EisTshB
THQXILoCj1/vmbB1qgDms06ax7Q/m5kcRQrZRWTVMVyL0H4mLNJSXXqLN4ED05gOD0m9PoP1QvGS
mDU1gGoXJIXvNv1oI1zXGZvOj/VfLhSJ36TtTDc+nW3U1QyWdeZp93rDnpFrdizZ2qNI/5gCsqq6
HkLtfkbHJHC1LkHi5uFt7Diy2Fhm62zMhZTeB93KH6+oaykYCpHlkw6DMOP/vX4he232Cp+dRnlw
OScaU4Uoa+v/zgxKktKjT9CSH5jtQ6hXGGJMtWjpIRO5kQohpS3R4b0bugLBnX1JWaj9d/Wi0+S6
DYsCWdJ+sBKy0ARYR5HuSgpzDfKOwCigx7Lb1IiiS2sUlsRRiMdrpsEUIMWLwoyacKZrUHhreMAW
z2FLgjBCHj71Q6+iz2YgaflCuX6oG/o32KC+FA7R3dr7rabwgBolykV9mqdGJe35ThkmdPbCffe1
e78j8OMwAWbU5fSBvbT3Au2QzVD6E23SqZvKb6gr4yrT5gkZh1PJgjh0jp3oaxJulHRGRhyYHUye
OeG4hTbNck/JHIRPr91u+vuHstQUt9bnW5ju9Xqcg5eR1aTifu31eWCOZ9h1ccZVSmjfZhlMWVNi
Ojn/MeoQ/FLDWSL+HV6ryLOqRm1e4lgrJItg3MZIDkYq5Ss1RwT354206/NNF4pkE2+j5mr7H/Kq
4Va2UWDXZ1uHqihLax54xz6LlZMqSLkv24ooTkzqgoZvyr9t1na+7d9nMFS1zquwy2IFcHlmudce
ZahMp5ENKarn/5C8mLKFckaM/jLAd4WsuBbohMJkdWECsYhA2yPC+YAdcZCx63DgkAY3XdOZ3GvG
TLbpDCbXdBlRXGeZmWOUiWjd5IUCxh4gelIhM4xo6tvupyhHKKJwORN5cofp0IFawTVZk4X9BDme
TKyythgAFIKpaZi6WT5rVHnO+FjwOR52H5Re32Vdgs0XrYf7h6c/7BJXIpBscbK24QOWZX+1cGhu
+Wqbe+ndK4ZLeR54srs6/gEMOTR/uVPepu6ePP5qclRHUmaPNS9O9p/vp1gKNg6u/T/pf8bRx3x3
1zYiOxyXwtwFHbbbLpvA9v07AdjpRB9sfoDxbulNCTwEyBAJjnPTn3rwj2PreiefhKpUbQUoQjIg
o7V3OlvlhGlZyevSf1pmObu7t2UABnyaSLMYKDC6xVlXeP918ba6yPWQcNRXow3XWUgwLeY5f+QD
WpiOl4lCXrulvDVZ6cn7FnIwz8HEM8F6NaWD4OyyA1uHR+ek9OVjruqczKJO9mvlfxxv+sImTT7a
pVolGDXt2EG+ssQEfXidCEugGdLUZsCGINY/RfKBapZz+ySSTut/trT3qy7HiIOgH4Q+VtxvyJo6
tvSVNmlMJpn4fKStzHaXflXH+/0Cy3XQUN0rnwwFEYimcKyGz8hIaHqoO3NNKlGBiP17iqFLpmP9
QQXO+CgqV57u9K+IJnKiXKbNSjVPp1QSJPyKwfFLvZqozHaJKS9s6tgxWiPoIkXOUjuztjt2cyNl
1VPjqLvWmhLFDU5CauDMLLndAATavBPUaVyUpas8aV0S5+6Rtw3TtJCUeusenMBGPrPYKYGjflAA
w0MLLHSnDEbVwTAfCvzgfkiG0p1hM9HO3l1CTa/FrlIxnWRcJME37brFV8GOdb9Y/oAtUppzBHNv
nMaBdVcEwAaXwLNKk2NPy+zYLhFCqZDCQpgKRXrGgONk5N9Kt7/slRggZvlfjl6/QdVBY/YsckjE
CiIXjJ3NUt7FuvH+JciTPq0QhZVs84vd4yN6iW29VwPEwJ0JDtBMom5M7OYG/3xvgHocbAPshQF8
mBTmDDueZPOl9r2vb5OcmPEWxDa7uug93qHxTobhV8slO1jsDcGPLn2goVjNrb8z6GJzVF3E3Z/m
H8ULJI7/3dS7g2PvJlS5nzTUBP2n09C/DSSmS3ZbwKzWdGyXNNo3Xk2/aOmXh+RSc6NsFfZePd4M
C4tZsG7H7oAli3TE56ZaeZqvXEKE6NeCOyqTBSXQ1ssOjPCPDzCjZ6CinivW/J88o25rQFUQ7RU/
nYabJJ5XNOzccgu5D4RigMhHmfW+vSrJN/fqczfbdmqtYb44LSDlL8pZ4kVthfj0RaCfOkMtIEoy
mPO657wtldAHNV+yqGr/NzVaWQ1lgldCiy2f4ITKRCxaaWvaoVrdOXqxsdn5p4BmDJvjeGbSPGlT
SnE40Xw3aoN7ZUa84D5dAmlGofq3Hr0jgi8dXm3V9/2mKdegmqJ77pYMu3ZKs2M8RV34fdHNKCGR
ykGOHJPW+BxQBTTqUawyiX+kaUYlzGgJ9Yg1oqyQgJxEozm2l05+24mGf3Uqooo/nuf92tLNYzxA
yMBKw86qgKuFDu8Uk3I5zRIoR85bla63rvguPFbVksXXy92THEPg80kNVvZsiVFm5xKeIx3NaN3Y
wBdHYsAyJhQf0KHYnNd6/BWcQ3ZFMqhUxysxE3AOTBJJ0Y3Zxsy4OjUe6PGr0y4JzB26YsqlxjPu
FQmeRQ6HENufGLYQK5oW1VUau255SNJH+Ty4Tn1QQKeuG47uwky3ZOZgPUj7iat7EtKNTVaZvnQj
CnLjeAJNKWwRMWiztwZr12AbVSaXIgseOb5jMVR65HnhrqLcpZTgqCm5mkXuuYg1bAzT/46hU+dj
ahjNMQpcy3pBeftIyO7F7jkWYECurEXn1VK+yK30iRRtXdxuhKESGVSy45eqROjYwh5fBUQomT2V
8jgZPKj/Uyzcrs2QDibn5cs8tq0+daFX/FY+goqg+2j0kR6yQSmde2tX3rRxRurShU/igEr+fNXQ
MQRjJJywAYQLzlY04dZNNRv2VOPwtlf1FsPlVeH8qNAaoRxJXc5NAt2nksmDPLTnN11a4NNjxYSP
+NyQprtAFr1cCOo+V/XRTWI/e08zLD+mgB9zW4q4fhJ6Z/zppvPjhaV5YTsN+SWDRlc+niCoIhMN
MVnCgBvGS0eo4/ig46KTwY4sr7A7qPls9gGR5KJcIYpWK+OKIftVhdQwKE8Wn5CDDNrxl7pRMyI7
4JgtAg55c7fsX7T+WwqYiTxOHMwweb+dDoP+YkYaAY5B2eXn1U7ORGvqnNnWCTeNYlDALFLq4vm8
TdQ6uhfJf3wxot6VJdepEwyJ0R5jvHmyqXaQX7IUw09sT3X9b3LWo7rcr8Plg6ViLt1LlGqnvz30
8mcF95vaJG4FAcjOR/wwQ0VJDEoeSOOb1q5UTnVw+wbBR+8XwUN52Q5Nx9JAKZ/ERFxbuuDYJb2f
mjwyMZGWQJxa8VjGozEMz/GojvSGk5CJnVcgnz+8A0FhTVSFZlgYxQdfy6vztQ5KpAFdmNxwpEP7
aGTVKY0sxE91kpa+/4m9vlc4WiFFCN6GOFH3V1vjW2rzDllXuNcILdxAipgsmwndtb+urB9TujsH
guDk4f43SlA7DCmYpsMJb0I0Ro4kHffsZcfHdkEYU2BoBrJRUdw0Oj3sZfXpJFwTF5tVos3VWiYa
vTWQMMBYGQZMAcIlb4GNISINYeEMJcQC/HKOfxebE9NVJFDydJIhwyeFgzvmUlGLDNIWq1HLEsRc
A5V4JYx+MyDGy7b5SP9dGpNAfGq4NwdEJ0M8to4heUo20OScONJ2X0iVqy9GxFNHcF8ZeB1MqwSU
A+gSl2Kg4Su1jsaBh/VsjyprFmlsv9FSq96tQgqIrZLMthZOQ418zy922hINeJXvZNwDLUYeR1qI
bR2O1sHtsLe5K6cXpzZJ+Rnk3ovQxBRgI7tpDX1gbJXX3YYtf82v9aDGJMDjak1WgmLcfOe3Rjny
y8f2ejk5zSs7vhN95SopwtxI912nAPTFaxxRFhmKFTOrnAy9NWKAbRzgFhEUaL2BMHBY72Ev2Gj+
8e/U0Ax6Zh0c901soKbsB7n3F0VD7tfEINdRW63Rhf52ALRT/mJZHZvPokwLjSEkGTYfcVDjl+4p
glHOJJOzydvLUMK+gSIw3yUhz6VworafQqHLSmhomASXXK7CwsOhnF/hBW0QGhuJcDNmhxLyVpvt
3BvUbGgl4KLsbFxfV0bh4/mdZxjqrbW1ijGBDU4ajIcJdY5N2tJDkieIrnIcDy/H11ne/hROTXeS
T6H3hdRkB50douFoX1aOzOHYXDVbMve8Kuhb+lFOy3vcOSvqlxN3Cx3korjjVJMWa7tRLlUPDGK4
YsKw8j5ZHaBMLpw+M+o1XBfNhOSl2eJgAGgMtRtaC9zYYPiBAej8zCucsq+ZCIgeJYdDJ69WoLVz
XFaGa/OVRjj2o2tQoK52dchCqiq1C+e4Zha1uP396KC9t2jKFQIIiOq1YO0Cftlt5VtQQVrtA0NS
qWXUS1zFyPxt6kbOqcdK5fiqOMReWF0IXZLrqN1/kDnrH4lM6w4yUt/Lypnk2vf+516awOtsJ7Fg
KK1Q368UK73gs3OJePStvf8qXXtE0RndmgMY05rUmpFQUgDC4CJDpO3R9Q/rhgXAuhibpyksCbeg
li3MbfDJWogxh7yiyLQ4m9SI9brJuRd3IvNDBTZXhRSqvo/+nFwKbsrOfh5glvQqZboua1aWp90r
XAm8ErQOeclUii9QcukJeJkdDeDUHMuu92RcMw25htnjXmlg3q0kI9i9TGHG5+e0uIz6aOPEl3ML
lmYeRo2aAILgDpptxpfk9YyHFcVvDIYDuU+NyQP4/GAvu0luNl32XeWRfIidhzhg70LIlbAVpR7S
msdJYXcgxclahtfoZadUyFlOHow/GrtP/H4bkLymQJENeHDkvjjFCZ6zZOw2CW62WNv5XapjyYuu
MlhNx9Q1uxIwJHTYK3cmdmVocuDQM+JPdSEwjGPV9FhSai8QQdruBRy9dvxiEd/ptboyLZKhM1z+
RoUrGJ9TYaXdX3Tekl6CtxvD2V29LczPruL4eTfxFZQl9hcB6Z2tZyVXjvtD6lz21VmeznRbS0GE
0MmXonESwVePsH3Vxtf9uMd+GHqTTiaJDdp3W9fT76eNmA0Bj7nm6/q7/t2PVm2v0tbHhDGGBry8
PCiicz0h0hdJgQ7BSVhXCLBXi7wcWm2bTGSLT5lK9s3fbKYEyyGnueTxTFqSJZPuXs/pH1RYFE5Y
O0JIauv77soexWvpDoluJCUuXAuIgEo+Xuokuq0JP3GLebm4IaHmglWLqlBx4fv1v1suiq9g2Y9A
ws7hx+uosWhRMbW8FFI2AuhpPML0tS8f0pQlE0gns9tq2uJDXEgGF9ShIVrzW6Ct2UPABxgVfgLv
120jpX57kE74ixBcoH5SslKFaf8AQk86QujMkCsyPmLEBEmvJi+IUxgg/ll/80qc4NOoiA/T9Ihg
EAzIPhNtIC6KpomxESvSDs4X3N3XgEsH57hORJZWOm64Lc1bMo+pWtl/VCoX+iY7rIiwOali/KVj
okeJcB+MmGUeZJHduEFTS+lAqHQ7/79xctXb+5w4aIb6w0aiPEcesQd5cwt7gYAh1y1WA84GGUpQ
sdO56YsbXJkM5dPgouGB2u2simpahjmrK9fwXA28fCwaMic/cP1QXMx1taFVZGUyFxWQF2PlydS8
4pv/Fp3SLQDdbug3oNWnW3MJK3qlh9FqxpJsXSgpAgPkzSH7VQ9VU5AwTchvaGBCJOd+v6+a5ssv
8WZ/yzCquoMFLcGVv3gYak+bn+raKI+MFQVaux1OSPEP0Gn6SCe6swUJODHESAPjj9yMpow3Ubij
l2s85wAlPhhfKEf9jbfMc1x83x7b9UHxvUqVqsWRNwOyutzZ1r2QCuLwboo3Tpnmi4N2SZzeZa9E
RnWWXZuikvBtk5INwXFh7TaTB5emrfs3TgUiQriWufOazp5JyY5Oy8gjr1K1Q4ICSl3g9IFFrvNC
/dblv+fii8vD50jysS4EP3x41xFR4925tmNPw/V0x2I6FyMUsRh/6ZP5b24+flPxjbYfDZA3MJzg
kkl946Zo5EUxrR+Mq6WAGhxwmbgCJm6Ee9CY5Ms+UVZS9QpZ8fwSxmdMJJJqPd7xq2GU45JrT89y
rdjdwcDxVYE7KfedaU5wZW/4MBjFbEnMA/eShK5NGL78kjxvvdIKb+B4lY+4jW0q5pvfoFDBKmSS
1I1jxj6G9QA4LWcOGWVQ0n1/ex5P9xOALD93FWjh0zMTN+hNdCw+3/JI2xScGU645T9iBIQEySEJ
xbJoM0BNaNr16BJ3vmzDHPslrXDh45ibsS/216e/og1kC5AH6575JDa+rju0DcjajeBMp9leg/c0
0IlCGHXN+g2CH/qXayPJ6+lthzm/DxykmaPam5qeyldmiv3GYpHM4khm8d/TcYim+fLxjL58entJ
j1c6LoXas4eS8QOzj7AL+eLFRx7YbABHA2jGUawKjqWwvoAeMz8C0TgdxYYLgf23ylue/Pk/LksI
UrcCZ7QTSsHcX2jyQxs22rsey2KrRClxBuxF0dtkn1m6BG8f3jyRJ+17EzzymHod05NDzphiAS5a
gGZMOtYSbAmG6U9GpaPwr0qNraz+66E91QqLjBA/27LQuZUD/afyGcEmwzDyic70GmmfJ5PxU0Gl
XY17X8234BI65Hk/ko9SaR9Jw5/DAzU7/BRiUUmprCsraInw/xosVuMDsuY5KTMQx66+1aVwwZm2
W5ozKHuXJyMSB0DWqW4+SDqp+ZGPlMbmJ4Fy55shxNcsEejxsaAleeCGILPZiYEdJhUytalN84B+
56CIGC9Uk/+oO4i5fbZN2FRv5WaZxpBx8/+NAj8jcstbFkrbTXVFyQ+dlZctf5iavN4p7Chmt0Cw
J9V9ejiOlxm5ENnR3mhFJYq7nkjNkKUzHQW/p/yMYKTdkUy/bNMazoMfNjRWylJA3fhtXWUFZsXR
Vv6FWG5J2/+C23n42fDqztOCCmJ96T2mVTEYJgTHOswC4HzoJmpN+3XzGZkh5IN8pDZ74+PvegAL
XfR3ElOjQ8neeEuSGSiZ2av1c2fftKIz5hRmqG9c3QVYkNWzbSvTYOmvwW7voreTKrc9ndoATmXE
G9WILN9GmaFMevLzJzYW147RELTziiry9/JSmufU8TxmPVWl9DiCKyU0yFmYOsTiMp9Ro3C6oBmC
8aIlZ/7jS3aXJRuS2ijXadZC6fk2n+5IzGojTPHKYlQTiAWgQl0+b161c+PiNFFpAlbN5QeVYR6Y
MD1I9b+YS0cJjwy5upWU6xIrSudO5LIIUfodKWX58+eYlzhyPhQntpBN9xk0I0B6F7CWZ3aA1G4/
HLUkN2jrUlul9MJcjOw1XUjzXethxc8p3UgLXiLv5qy3tZtgTnrmBIcsctswY8zcGC2HM/XdJtqZ
h2GxXjH7EzLtrWk+1wcw5ie7GdIJCI/hxV8DeWgmlw4S1ZKOmqEFhNuceTTbi/Jks//lS3bb29NQ
S55ABilOQGrfF1yS2ncZrf/9m+dnm1sjsSLkc04f1wgUFnn3byEK464DscS6m5u7iG0zRLYuARAE
yP+3aqGHvSHAQLIQIJC6b8I6uMbG/uKxQZ6YBLmadmRvGtsW1kAYVMEIqMuQdY3ixiN4CJTlDc8I
iOOWumAG/5ZkVqV50stoR3st9cMET0xIeJd/LN1yg8LPdt3ebxUlLAY8sqsm+fAE+RSzcvUUGprD
9MTO+KFNd6EjajuBaT7qZFcqdOiQ4TbBFhw1pWKfAE3gULF8NZSRSrGysMZj/QQjYn6fTGY94FaC
MIWm34gSkOtwiq6Gm+w5nTr0G2npq49IqezJksTzZXlHATJgpYUPyAIcpPqpOR8CveyHQSuKFYXT
X1itWMChQzIm/upo/cHyH0Pkw4/rdEuunOEHo10nsN9INTTVjyrzwVLg/wm21q+rIm7i2gy4/KlA
OYFT8cloQseUgRpunu8oFmTHNsOqcODsDM2xT07+1YnNEdLwZakuz0R07vgBomr1C3CiGNNrJTe5
a7kZUV7DRQuFbJUNcmmSePgOLU8vuCm92CjQkNm1kn2OTv7BYWhvKX0QtyQ2BpXzV8Zyvpq+Jf5H
J2sdHdzEYxOp/RTMT1GAwTtkZLKCm/rmC8En8mZviXcS8Vj2zQamGSWgQA8jvpRjz0/bKpYDRT7r
o+/DwmSb4kvUeORWrQvhHt9eRFnuTq4JdAzZKmnQok68CGHNurfnLSRYA4emdHCAObCdNaPSkxTv
uo27sxINSqctFp5nksoOcCMGiCd6103nGwH8fGdnu957p9KXBjcM4etNrXPkW+nyL2NSviE8vDDF
uD0n7yWxClkQjIZFAiqE7g/spGapw/i/WSvbZcg/xQro2dlAujI86x5pmlqtqzScdEIgjC1Hcdzy
+YZuQOSeJSx94AqdFzrETwBaAoeQC0O4oSGAW+fnFJLSNsTe5DEon0cmR42xkHK6xDJLszkYzXyd
Q4TnpgfVUjTa4VLTIHHNVgRkD+wzcutR8cDUEPIixHgAfhl3pIYhBT6gnn8Vi3+EP3l901+NLlHa
u5rbuDFB0QTszc4QksMOwixNZAJHYI9ynFcyWBMNlK0wmeKVNNYIkS6+URoNbcUDAFR3S7nOBfrx
dq0QATd+cKX60q/AWXYiXmLYF7+DBTI2rTBxgJTYgZhF77BjUJue0y0M+SAYxoIXdPTGYuoh5sE/
FyVK3LE0OSUVhiDqGqv781aqlYf3USOzgq/res6EK8hA++qz5ODlv9bsJVPAylxY13xV8THqATWJ
tOkVtfP6AUnvxzuBn+u1rlq9Bn35/t3+SJvJD9zt1TeErb+l6djxcmTWybEdjkGyGkw4zi10obZh
kZzcax8bL630x1sr3+WtBzirfljXK+GjNYF0BwvZfK8oGBYjFt/2oy2BqedUzr8J8hdwFpqfXcyd
PV+LB+BNu7MVu08NkuVIxU/PSjJr4Lhgc4AGdaAHx4MjGIz9eKWop3IcHMbkl3TzpAkhjkvnOYx0
NC6uN5wGIQwKTaJkha+Eo3h4VwQFuEyibJmQ8EwnruT2WOKsZulqgFnCbEMoKw8KgEjQAdW+EwZr
QG2B9beVFXxlAku7iiwt0Pl24u7ojAI4FQlurQHzdGttDKaasoGhoZUZCAZcQFdbG0dzXGv/MN5r
J6HHBldvvY3TnzgiSv/a5RAGhTrj08VBsxM9hxkUvxiHPcbUXDPU5c6UCoHPTQDu4VdUNQCNzOF2
Kc/2pwtDg8wd3UTz40LhBUsmlNuKeUBCnF4mqroPRSJ1K9bBfdI/+TNtMYQhpawJ4F5yEOoJ7re9
weUfRrBtFhxoKAcRruefmr5mPCDaR5qb/sH7XVtT+h8LdrDnKZS+AICc2VI26Md30wEsieGeugOK
GtvAxn+GQwZdackI8lvoTKypHKPDbrywfWX1SW34bFbjTWWA9zT8ya4EpXhsMKXYImr4B2FK7GHi
dQy7L7nkPhL+szm6jyUyRCLcFbU7ZcT0k7frr18yKPfDZx3Hu000NZhYf2hGZI4j0yKx4/x8URqw
xXPlPXCx6eeU9L5i5WkKybXigutwZ4di//D3xzdt0J9K73pySiaUn4yEDHbqXVrtkEdXOVE7jZwu
M6OU/sogN9mRdObEJrUReexs1mc7yAEQKPPKzfEMbnJ/ar6gRnw486thOyykuypBF7tu8Uruw/P6
8Gy20w+46I/872g96889Zsl8zY2adVGA9wlJu7ZxMxTZlJBmW48dLOy9QHH+wLgEQE2kFHZA0sxW
Pls0zSA6qeZT89pKviXI4sMj9m0irt9Nw4Sl3Z/Sf15RE5DWO0OIaipi+LwyQYG30EXRpnmwYS5r
MRNogFq8MHJsvkN1brjXLweWSzL/XyfsGoZnvnIbEB7cAYszlbVP/xSeGe4Qi1VFxK6tBg1jvHfz
Rk84qm0NVygwSN6++fbgyI/weLn/dB9JYyhJ2qLTDootqP6RkjHzI8DaWQ4AJv7Jwc8q+x81msjf
PnVCaJinB1RpLZYJ05tryacLSVMrzRDcIkHP3kuFHYq+ZuljwcbWcEEPBiK80V5pUahUSyn5C2uX
r8oiaqVZdQQs7j+WmrvO2HnXEIg/SE3d56m2D637/xR2RInp4R1yt+xcwuDAw+p+l+yQcWVKGTPN
uUrTRa7VsB5YZ6xpo/CsX55pf/MxzV7HVcQpRM5Xish5db3nLnEo677C8UrPWlPp+ErbHhjkp4Dv
2vw6GC7eRii/SKR/V0ca7NOvtlU/5b4avGDpxjYBG7QkQJtpNP7jS3UKqYrFvUoOZDO5xJ1WdD8i
5iCzJaiDhupnTunt6xRBattmNXvFLBXr1qJjjdbjDvrt1Jkrxe+a07c8up8CMtO8zh3e5DdPmsDc
YQNPjvSUmzXl4X+imq7OxXr342L6fBczLbMEUvJ+l0ympjSLWo3rYS1JX5G2ECiVR2m+mO5BJBa+
3SLd8ZX0RknNoT8H541LsJ0Tt5uHx4RBRYy3e8KjBf8sNuWSH9fJwOsYOtbhCGKY5H/LHjDPUwbn
Qq3xBsbolO4FijxY04GTGAVd8xzgW4/DfaIBHJHoQ+FHUYgSQDcB6Fb/ubVQslSE7BpxbqivTWl9
LunnEs97KQLYhNcyeP5546kTE84awEHEcERSy/QL/9PJvCbIQL54agVOMhxjP1nk5vr2eqPLJ8BX
mnv29tm0kNAIY/dSOhuoo9zhApF4TjqLFg1Vk5WCkvgChAOplW3osNXJgr8RpEQWABfU3S4LPlad
SAFRTkgYLLAO4tIwRnan5eRUogk8MOH7uSS0+DP32WEBuiH5OcL7awTElGV9L2fyL0X4b4pfK1Ce
oqR1bCRH7+KzHp8fzjNRevibpl+47/4wn5KPf8rGzIjzmJKl9a5Jx32cMm+FYkYBlwYbg3pZyxBd
cP6EX2Zpco/ipz6FuCidag8Mtt+Dqm+cc10YuvjdFgNtiGUGL0KILbkKuFiu5+nQ5aL0cxa7w3md
IUGZixIniLy3mH38HpDyH14/+WSL7ndSYg6VpwxuW4e3wi9Uk8y3knzYzckBDDoRum30kZecPWXk
Z7M5wLDOh7riRj/GrkeReXeNBLTK5MiDHSP3aHIjBYXFt3qZRZGDGJFFnwjf6tU4JZS7hxnn45zJ
5EP40fy39/Q+Q1L9PWQa2r86HVSoHv/ubrd8Jfy6+Y5xbER7FnUknIeLsSfqcx1opMq5INUAsmzy
cdLnkOchBWbiOvFFvqFf/J2pj/xVnqHcZu1g6ZpOrlKASbr7gXt0lLFQ+g0k3QLarZiJaMWuLlI5
qaeK/0XSltpjgziHykC/W7c94v11XLnQaViB3S1RWdI+7op+oCRU4q17vGwm/nT1sOxjZlVH+O66
dghr78gDavlxO03ZMFmvx7Qairjeh5FEgTQ9c1Pp/pYBqYRF2qUN9N332l8+Kb4melADnxPdaXPM
g5SOI2v6AAYr7DNS9PP2fEIjWUc617HDK5U7etlveyhKl9hfU2DCYiQQZFQ8w6+LTuhFeTDbfsLV
sY3YeZBYXbrPBBtjMUrn16HF9p7TvOQIR0qNVZe0OdfQYVjkSGKAR8sBbWT84tNsfgmZ1UXOCc6d
tVzyMw4Bfw/1hyuwJNYBt1hpDk3OporW0u6otvY/N83BRiIgCcC78ruaXS0Cjf1OUzaUokqdXxTN
dqolmO99FpCsUw0e/rWWaFccpVzJ35CHcgHgxxGXA2J/JUf4T1xbE4A1KeV29ALo6Mn/8wS1fv/P
vrSvW8cM5BWaHpZ9QvOSFYZ/FUcpIDkrHpKRTnS+hLcWn+87D6YTzceb8j+Sp/Tny28Mz1en76Ri
oPH+quTT5lKZPHrWMIOy8pO750GiYrlBW05mXtovCqxoEoK7heIKG+/0I8L92u9GoTPY+Z2n4AZO
YB5a/UuFvY+lrTzWvYYmqn11prRzL5gjLAfS391NAZQoZ0HKa0rq4k5zftjEcwFqTyzGD4w2vlMj
9fjV3/L1Lfk8Vab73/sU0pmy6vbiwjRozaiRy1wtfpvpVHBASi2X/qFlLPYhcz/fc+ZArHBWdwvd
pPWOlG49xYK24DSiZdIQ2PBUN7dBfyemb709lJgJcNnDMvb/MZCdsWqX9XgGJj/azwIlk0kB1sLF
UF1/GCU7wlcgpEHJiTSszh8Y+yb9v7q/GuHltQpPZiPF0P5j+Wh6Op1/bulTfK76RAzOaXMNFjaI
Rs/hsEWv921N2hGmz0/paOpbP7vBLak0+DTvEyk0BGTytV/bdpeE4m5hubeAtHb+WcyvM3xtM20W
pAhoJ22rYzPjvgo4/p6ZX92E9YEjl0VCFygk70Y0p+jvqLiERB/NLDS1Y2mSK9QzxC9NLEQnE40W
OBz4LD/BSBE8yTON7NpHz5Sazy1yR75Iu1ox+y7bRQAsrvO5MUwzEL/XIjLb8w8ZVX+ZA1QDJcAD
ny2Fiv1NvfMcAdUOGm7jkTPTiLAQV4VMWE115/9Y+vwaNdfeeWY9k0skodz9Aj6/AEgcgPtvQubJ
dPuhb95A/i874LoaMACTN+drRZS+jwsS7k+6jiVGwU2FUX4EkeGxHUyLfAB8RcVGMg7o7BiOh+lT
EKcCZCdv84gKrfb3RYSuT4Q5CeXr0v1FN/QSjgdvwADlXLVALJWY033yq+tFOyXJ3d3TBHRHOzaq
gdTMi+D7oOesODm1RnLV5bNNK+oSlU+1B4aU6nkzeXws5YMDTfQGd98idilVSJEzAVoc2IT/oCqs
yMtnj6CDhvAwbZeQGSmXq5jejuCWrRLMowbzGRdFgS3zH6srO4gx4EONwYIZX4Zl7uMm5e9OFHzf
s1IQBLjzKjbVNI5btyTNAcsSa2468FWErvu4RUiPMg6MvuZkIpTLuGjv1R3Zl7zy2jYngW6yeii9
NfoX5EK6fXhq0+WjF6dsg9UF70hNRAG9pyNMb9/+JACCT1l1j032c+yXSofyGpE7CJNAw41HGGES
obWQ72RdEizbocG2x4ESYblYIPRHVsqEnoE1+9hnlrP/0oJUnyIx8C2Cx7WBUVjxZ+AOGe+gspsx
qh9XEoWp6WaDgqpWZKZbAeWg8AQbz0A/m6Y7DZEXZUUHmhNAw/ykW7Mg06oLBHM8CFt4Qh9oMlje
taNM6IWHPy0y2epY2vofqSjaIRF8hpmVYavV5XLlNHsjSXgXV+xkGdSmfr9ArDI6C28oOnlM186P
i2+hSrR6unHz/ycTQAuaNPK5yDNvKjzUr7zzOjFYcX1wicPfqIfi7q0kcp9XiXsB+V9bu4DmDKmT
sf/NAJkDqPwKDOBnQvyD85ji3DkJskSSiInTfV1nHl1nFjL81bc7dJd4Tn4HOSwm6PyhOv4nal9c
MP1f7wFb/L+zb+k4oPL5SIeKwpPQCFkVVCgMNshdI+01jszvcL2alTVLOL6AYm4ApgjTGF+nWx8j
fyppbsoVKZfjvkeZAW2IsLnnTeu9DNPrDjSvcF0A+dU4y8ikP65x4Yp0hCmwuVwOEE/OjlSTbetP
cHSShg6GDC90dOieWDaBK+Fqsix3ou1nBSO9vqFhlEssoK0KHtLxLhuc7ZqqVXJ0kcB1VQHdz9EZ
PMBhR50B3QrHbkV6G2q/0+508vN01+fIKhFKi7bg1mbfGUZvj2ddUYB924+ma2ptykp77FW0kfCn
5N5UW4/k4N9JgqP4jIYfzbcRbU9PkBUkpkH3O5Jm//jjsNM1qaNkrQQ6vxog02meFkp5T3aPjXdh
xD06p/EPY3UraRKn86JfDPTrLy9BXldIcW5HHyTelVY8Nv+YutjPdCZqT4nNgoqjAoKffO07Wnjs
/WYQc0HqdlHnvBaM5G6NQ7I4LfdWuFHi0nklxO3jFIzaGEzD0DcsfVGUKBFddjsCYQmt9asi2/Sa
OnOtVIWh0XugpigTv3jG4k8bdLXIU6xYQqwpHj1+3AIk/cJjossgCM75t6acg14ppgSl5hhNvBA3
HWW7sx8CZnz3ZsuWYxmwTmsv+OajusX/JZbSsTlR+w/7TsQpyP84puIF3sVzxTl3tQKhujxrA6PU
KOV/+Q5QYYNj0F9D/0dF28a3QtIaXGvoAbw279QGhSjDNfnGMF00DmPkpbP3T46vz6f7zsxOlAme
my9RYCIRMaCFPgAYAVeXj/HTudy8qjjD4hIvNYMat+lS/hJ9A/tTM0yCpU+CWc6Wuh0VgL5wjpB8
scGUBqF2INhoBaYemQZxrP+gK6rxYXu5XX2mPhfBSc13v2Yb2LJIVi1bE4nrPXURnCmbfA4GhvCb
tegEAtVWUcPL3Ep7pn6w2mjDRxwYR9ux0YlEw3n5iFgl507vimfDVBOjdoT/x4F45a0jGFj3fIFs
svGQtE8t8OvW+jvzSXJqgyfgzlP4KTxN2aqTYXKea0JB/c7x/AKShiqG32ijm3ZqmT0LPN3v9cYs
ieWz5LTZu2l9rWV+rqZcLsiJXxJu23vuy4BXu9UJ9KnNlMBGyFsdLJR51huJ2Z/M+siNPnbK3hST
MBnjNxt9F+cYZKm4WWdqihG3usIq+l0yQceBD0sYnE94Q5yje84Gya+h+wFgc7sABJd4hsoQcOSf
IvMG+LnRqKoht/SZelR0OkCEBp8CU3XlsPUhhT2K6WEQWv3Tm0VJcNMTlFlVlcMJ/mMEI1pCbGx1
8LqzPidtTEon4+4tC7Vtrb6tRQ7Nut94rDA1anzvf2NajvPSfAQ8WelSamX2VcUiVo4vPFmt0sSP
2kdBl2DNWgsbXeVP0XIHXKAX7VgHdoyrKdsNPnmcTBc2VXUqrfnAG1aZFLAXWIwTkq8SLlElaq40
LPcIlD/oxUYTyvk9hUDthImprafzrrnkGiLi7gkR/LjbnPRt4eJnXXSyE2Rw3tubFniSgvGNkHZx
OxpmW1VwZsLQ9i3RJqeBgNM/BIxVg1zikfVrigSxx0Vyp4XbDlYQnXFydqWRD9Zy2rhki9fNFrxd
MU+ZcbdeV45U3aoyMrMD6mQTjHK5CT1/ZA2H4+XU5UZ/VmRuG72WKbDBqASfbaRmtZ87JkYD5tfA
EHllUD367H618cpg22Jy5lmqaWbQexj/eJILtdxWQQKnKgthSWmUFIZm1f5nkrCgxykFBN1CLm78
zKFJ+PaFYIvL7ah78kNGCnQQx7kaTQAdgA+FbA7NwceHZ2ltf9eL1bOPVFt5yo64oJvO8ru0zO6t
QQPL2PcXfM5Zbp7YGP2NE+GTvlDO/1V/yqQopOCkqUojvQyWw62pYy/0y4PgAqfJppfv1erCSMsE
WW5H7tNNaV5PByQ+oj91IH5+eZu/oPphrF1f5DDKFvW7Hg6fnT8K59Dc25XXDXucMWlFpiTnauR/
G2FTKbSRr1ibdKw55n6rVNgQg24vQhCEhzcQj2A73ua5L0ZBWP8vyn+HFmz1odFi57a7A6er9IRC
THx27wpaFuiHPlI3Ryk/ZAkkBHF9LxgSm7YfQIk5HdR2Vf5jhoFSOmSWr5erKntfurSkDtrybsdu
RRfuelY5MtEkZ1kDz5hRvMeMq0YjGAfpRyBSIwTsE3zwpxqjY8Ppzg50KpBRsuUdzINdGRb9SwM0
2u4e8VlBvVRSWl018Qt5wyva+7JLMcdDe940ia2/8v6W2Fk8MthyCsZj/GPWt46MM3DzqPT3hIIO
B50pxgZU4JzHC2ZpeS3UNGX8HgtypHx6foFKpR/V/VniqOVXbBHbv8VD/QiTQ9ac+dqhTLULl35X
W+nfyLA/r3CgWYQHBczYJGu/Vs6qF2THZ9b3HfZZFjt1YuPCtKMomlNYDcgScRLms7apHKNwvEzI
m3+vd/K2NNLa6uY6mnbAM3Gb8P42LJbgl92Wcxql1EYZqr2ldkfv/S6MaoLHYxZBMBMrpN973SdG
TOQN67guJp3spnhpNmt1NywwcoLhnopKt5OIze1aZm6KpFWOTiXq7rHKrhaH7nML+N4SzMkch7I0
GM3nfVFc7eENPjfdLzx9P2jhK43+fR5aMp9ZWFcN8OR3Op6pD8GaLUqjPjuATV0lYPCtedyOPl4u
mer27YtZ5goK3AXsPY6ZQl/7OL/R6czqV58bDl2ghcuZO7A4o9jY0MMYNP5qutH9OC0XjMDIo0C7
M5eVPQJOXClCwE35a5iIX9ZUuglWl8AUD7NGboQNJonDjdvV9PgNCDbqcsuIii78bFSocJ8ziPZz
8+Avd9L1E/bHbBbJbQa230Ng4fJcN5gUYrSpk8VXBc8tKRLBIeGl3FiVpmE9kAMsNzUfl1UljBar
y4hqMBFWd3zJvlKU9SKM0WlzH/syK8Y3OQQhfLSULVDdIQJ9WNuCBgKttZ9+aYcAM5BmP08CMjK6
hXARMmT5mpPPdiI65YCXMZB8lf+an5VRUZNAe07p7LnlhYipouV0Fha67JFfwEFevMZYFwsbDofK
Nbqn2Laiu7lxfpvUrVXD2a0KjwBym6fWr7JuqN9E2bl9ZBL3QLa6qrq7jj4fihCB4TVGukFNJ0em
j0Gttz+RNMbDQHZTqtU2qngfgj6vjlHy3/irwnerprrZYkWaCVpMciA4BsQwCLKWnJo4F04C2rzn
vmWxiDOMULLylN+IrcEOv7a/4j+6aioOZo6vZy95e1Xdgio/9LuWjEaiivczQTKy2lkA01RH0JsW
QVuQBF9PpwcVyBH/0fryDFIzyZHOADzpydBd2x2EMn0kNg4axsBtm/+vbz2tIfnHASyKPfblAXak
nKQKKBv8vx8hr/C3YQcMJFnJ31P//u1lv2ODHjfCnDbHYj28FtX19m6cDQvv28S6Oes16gX4tyw3
J43v/yUHz2MDwAeAyXLRDv0zbVWRXNUnmZG6YskP10I8ZEg+44370O03S7lAenpHeTac914BX55W
VExC1i48i3//bif/jjhisfFv/xpfz7UNpHlnZmyFNT6IPqKPVuyxRkJSsV8ZQ0FxlvcZOv3VU406
H+W0E87rjWMe471P90mRZzlBMuriPDjQxKp00VHqbTH8SP0F1L02dDjPtbGtqZtBZ+9uSPEIjz/R
35tGKWkcRpTQFAfkDhAmbl2cmEBSk2GrZGcfxQfWoczG/rriGPvSxSVf7LoHdHIjzx2NY4n/055j
MNYXU3k4JBwhvi48ku6hCyN3uv7SKBcEqgt6Rbv5Uqr3aNg5/y6MbDh+yoTrQ7B1qEIcko1vK0x0
n10ZjGoMem8kwa5cdf6FNTsatMg6mCld4+mUVgpIP4LOGv9wmQBmZh988Qa2sBA940J15XixaAmR
7CCEMpEEGKINt9M+X5qRNv0kPtMxDumxv2291ddMQH7es1Gc/tmSvaSEGflydov0N/TqRnKWZXMD
r2VQ3gpRKL3O3OK9/FbEjxcm0hKe72f1wLOBpXQDC4easog8MqJZ9Y4CpwsgbvlYE9dJJL94iPzq
vn87xJUJ9xZEE107fjwQ9duKk2UlPXWXZxZUb5Fr2mmX0/4I9+vjICZPOmfhHhefn1ahWIQfXlz/
+piqed+Y8+TfgzlupD/Q0/cYA5IM4gWY2KJ3tP+bNRis/SuEIxhUJ2HuLIr1NWt9PBlngNHocY0j
evotrXJ5AxbcpONe7vznKsF7JYKggi1mIcriMqRa8+uZKVDGOnXpOYBJYrHQUVwgYExUzWk2xMCx
6f8zZ5KQjJLd9g/OoSafZEYByRQT1ucQgUjjIx0WjhJYpFJrKJizt7EPsukOcU1DMfmN4TQCIbND
HIGVmKTDlLhRlIGlHDP5H0Kk9w+wN8PQOl/ia/mPNiAvhV0MOjnaDtZ3htMa2lug3skCb7ZD1TAp
HDMwzByb8jIIkEJhyzs91h6A8CuvM6LAQzK+rarYqhwhp8LCLA8dxsDcN1u08bk9RVkaiTvKCCKx
1rAMTEKz0KSB+HuFBnaobdKLThExhNACvKk2zsn9z9Ob+JKSkWAW2WTTKKt7K4pmI+btg882Xj2o
osUFewL4/ONAI9Ui1SB17Pdv1i5zhkEI0zSn4bp5+j7/DtmERSjTheDb9G2yAkcLgFgJ7YxAVPpR
T/Gwp8unlSTByS23OsYeknd2o090uasyOKuLfj91pPC05mcP9Cph2CBPTaCUjqXxlaY9VUCzqHH3
LdhO3qOzgq2X+YPaWUrvjzFv1OXta07MUhE9EBMjw5j+ynbQy2uMJNiOyxQ394DIKmXhgORj3Zac
k7S00RdbhCcGsZiIrqBw6Nn0S64j75IO2GS+Qh/wu5yesC/T0Xx2IRE634rxdkcGbYP0jD8PYCHy
DGV5izKZXLvyJ4rDCy5L+AhnFmlXLtz+LCAD08+e3xvHgLR03Mt0gdm24bFGggaGCJ9+1TDyK0Kj
6XOgijpdu9v+xfM=
`protect end_protected
