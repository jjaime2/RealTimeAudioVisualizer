��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?����K����|q8&�1��RG�|
��ǐ�Y&����ͺ�ä�m+����ջє x@C3>�r���[�$�%��?y^�	�sR}="a�g����巛���}���G��t�8?
���ཻ?�9��P$fsq�;N�3�Òʓ�����zڟ�ŵ�j��In���L��xt����E�l��?��߾�Ϣ�.����3�d"�9Ɗ5"�����$SP8�|qFr���V��hr��|�w���Sd�O�I1F���k��ƞ�;��c��a�4��\�S��,�I�/�@�,�����me��5ِ�M��俵�Z��B�B�0����~b�x�Tv �.\(��%$o$:� �W��K����k~���1�r�{È�_���9�<������I該�a�#
��s�ŏr���v��wC��&�tM�1��E��B�:�Y^�oo��Ndf�K�>Y��L2���#J�"����vRa�v ��{AUY\���q��4�;	 �{E�3Z���	=F���U^t��s0����=
�=H��i��a/��D�g��E	�8�N	v�0����3�n5�Z>�f�v7v�A!6�5��Gl��%��B)v��J��O�~�~qEډ3�¬��Z���r��膀�Ry��^t����EC-��-�wa},�􆮟��C�Ȭ�~��zbY:�ز�r@?W���20ͳ�TL]W����'Ί?l�躡�����Q�sJ#Ö�@��j��)Q\�,��Y�&��%��t^��$_��_S�*¹֢��Iba���a��6�544+�暩�qJ�a!�>4��ymo6μ��w>�f��O�vܤ��2_PнC)�?�[Ԟ��(9C������٪Y��X�ն`�S��6������r�4�I~����=hP�q�M5�t&���P���P��L0jr�(������* G������6öW#��:�u0k�rM%`�Z~~o�\�%K^+��W�ꂫ��H�����M�##��B�)�4e���2*��G�~-8J��Ѿ�����*� b`�!j���j�s�xS��|�Yav���7#y��^�]%-3���N騠^\M�6/���\Tx�2+�x��hk"X�|��Ǆ��@��V2��HĻ���x?���\�O�5<p���+�g���;��K
�upl���-������}�������s�+����|��`�N<E�?����6ʂ�bЍmRoO�U��J=�#�7�giq�]4�럢�U|<���! T��12t	��O�����M)UVTL*�;�q�c��i�4>�z�Xst��(�>�q4~p�R��>���>xͽ���OKL�����^hy�y8FH_�D��F�/.�/�����D=V�. ����\jf*��J���<��0�q�!{<e��ϔ�XɎp�t�2�@�9��0�V��#�ǘ�ւT򺀥���Z8@��ό�g��pp���]p�/��K,�X)�I*,�j��Z^]7e��텰My뛽��ڽf���twY�ma/yֳ=䙌�q�Yg%�Z���Se���|`R�����M��]TVĒ�����u�u�b9Ijܸ-�~V��!��1`�1��*3#�Z�E�&7����9H_M	� �������߯�iN@�[�v�w���v����]НQͨeu��Z1ˏ,����wm.g�N��aAcq��tX��+h��!!TU��z����~j�q`�L��b������}�ۙs��u��l�D��Խ�	_�[3��e����L�GϷY��A�c�g��
;��Q�^k�D��Ȋz�#����ۀ���� ��w�=S��i�RD����c�z�&��Fȕѯ:�D&���+���c�:Bq����h�sb�j)c\���>8|�����o�f�$Ыz5b�؆ioo���Ҭ�o�d6�. \2_�J�Fa`�p�Oުj�D F��ɎN����阸�3�T��fu��sȼ�aG�/t�7Ӗ��p�	�r��r��!ު�{�)Ձ�G�@�׮h*2_{��	�"ĩ��Y�[��a�v�ޛ�V�0=���h��z�8�X���2�����X̒��)�y��Hb�������8F��O���/���`�����u��弢�U�.���'��E&k��]0F������+`����,y���Ubq��Z���i������� �C)]�4:]�vqj.��&ⷽރT{�+��~6��]4䖄�e�3�c!-�^m��Я���6���o�z	 J��8f7&�cZ_����b�Ǻ��,�g���z��C��C�k:͉���[�+�`Jd_��f�;���H�������i�
!��+2�����t�`��<P6/�#�"=ټO>�I���2V����bIԏ�<�SHs|���-�C�:���dw��k�W�ȱ����l�ƍ��M�G�P$c��H��
���غ�����ِd�XU�V���vY�W��z�Z��(���1�[h*�mk��
�Aa���Fo"�=g�XYZ�5a���I ׃ṣk�ʢ��XZ7'��`<��� �u���/��M�Bo��_c�.Sc��p�����9�6B?�VoI�w�~�a{����$���%4��<��&rT.��a��j@�Ve~���;�s��Ol�/
""8B�bnOF06���"Bٜ�oPٔr�����\/S7`�p羒�������ti9Q���T�}*f�o�,��9Fhp����]]��,M;
�����!�A�>��f��4	����qyA(<�~��/D'��r���腝ߞ��Yx�U�R��^J7�A��+(6�������Lmy
�`֎m�`"��yID��.~��H�BzkQa[@�+�4�7�L�<�6����?�����
(����[��3Q��C��M�_4���S �t�$�y���鐚��|�y����s.Z�����G�Rx�H'�Z(j�.[�xT�@�7Gu�#��m�����d$`������S���B�����9�����(y�Wom�n�����&�eT�x�g�^��t�u���g�D�~��q�/3���Bja��� �&��>"�5��'��d�i)�nRtp��]�9�$*t�Fz���p���p�=�y�	�2��m�W<qD�m����d��楑�AK?�&�����c���'�Z�9l���
���F���WLփ��L�4?���q(Pg�"o_����� ̧tf��F�j��3"+L۷B@ki�N��it�1G%tPtj,C�j�����A4�xۻ��$�>��o�*u�<�tJ/|���Ͳ~>�	V5�C��d���O�^���	o�ҏ^g�,�g�,���9Z�N�f���oO֡�#���]W����J!X��C��I����ύfbX)�B]D^l�^��ܦ!,c1��aT��Cș�
����IcQ�U�?8���\�(;��?�>�W����t�0�O!���V:VN�D"�IB�����d���hYQ�n,�BE�aI����S�\�R�3+��вwlسDY`��1�v �׋�3f���`�1�e�(K��G@�G~#����u.��AJ�R�qy5x%_f�K�V�E�]\)����y�(�OJ���2?�u�w�� ɇct�y_!�MDM��T0%J�!þ,jKe{ڞr8�É-R����"��M��h �� ��R�؁��0i���cf�?	*�d¦�x���ô1��BmvPZ.x�`}�2h#���\Ⱦ������L�f8`�gV}��Ջ�1��>3~��DL���T1��V��h�np�UJ���Ax#k� ��"c@�j��3A#$ʿn�_O֒̄Ѧ�]U���[�A1�J<}�P��}�P���7s�^�֞a�Pw��6�1���	
i�V�,�4�1���Y�3YA7�/�`W�LȚ6�JZVG��Y���������M�W���W�OtF6�Vsu,y^�������E�N�&����9��ߵ���R��_WQ6���?�H��.ș��+ｆ�N7��H�1��)�F�Wѳ`؉[	7e�c{Ѱ ����Ƨ/s��(�/�02 ���v�<P���9QDb'���]ؔu%*���d��G���)g�#`n�6aZ-��:�E� :��b�(��A��EҼ����]O��$�Y�|F�g
��1�o'5�!Y�i����a�����W π�E� p�2@(K�?�q��Yuo��<+��`tFjc[#�l�U|T�5���D��B�^��%�1�V�/�M��N_P^�����m�u�?6VG�����i��Q�L~-�q��.'�^K�DG��fsY"?Cc�ABz�g<Q�6�?S�� ����{gR���VM���n\�ے$z�]B�ڱ�]4�t���(($��@iU0D��`�`��9p)�=q)��m{	_�)�^��؎f���`�4����krR��r��m�1�5�b#��`�����͛{��c'��:|������ʒ�ȏ��$��O�׵)������V�z��<��*�y�T>߾��Eʑ؍� �
���j}U�/��C�����