-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zAQWOca4PZdwpyNYKzoBsuTBWWkZOFKmkroXBe/5oGeq0pPSIMU0zfTq3dyX23ndJWP8vJZzCN+r
K3byw+6EI5PV7fqNqk7jtsndBhEr1pRlUkyUhrPRxVC5WUJQc1IvgjvrBD/dS/fVThLqMLQVTU9e
lpK+t06CwnGGXtJWTEVCHYQEdoAyNuXPa7q+QJcb12ulxNu+40n+3T4w5qE/fHxbTZNa8o9+hv4Q
0TdobgEBxOQxipV1tsAl8/PUkH0oFIjMaLesegwEnCmDDb+d+uzvz4a/cs90cpug/P33nIMvvb9N
sukKDfD/lwbrSukC4VQJNQF2Bs7L4Bt5G9fqXQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14048)
`protect data_block
BPnOzyr13ppxoFWUTEY6oJvaT7Ma4XFi6wfczpmy0csYSEQZUcImUyMhEVRPgVRyWd6gG+8CQXy1
2P1arqP7omzskOHfm1NglOn62Y13hyaE+QWiAvd2PX61hfor2pHqLzP1OVHvH5N1ADmvzh+YzRGd
1V/82zrrNkOa1jgCIJ6dVenj8oHw3WphdbgKI/jeXtW6y4wPrm3rydqaQ3Ef61qU6ZG5p0ckVd9z
TUdNN8Vp3aVlsDm5YMAX5oA847oVRpi0K9EUIO9ZDMuT1y5UPz1xfjLeS02HySmbOk33EbYPb+tE
P8SeKD83/Yqkkx00xELmYIGbSDGQgMLvxyClKTSjXrnjmeWMFVwKilLJJ3xnfzL+jXqDOiZ5PNXM
vFHXPHk6xXnm0/AxQRadYTFgC9K8t2zUlruyhvQuqch6sMhW8pawax3z66WPb5X81pmjELB0iYmv
DkHxc/jfHNVbMzqnD6IstHf9V0ktxnI3NiBM81vux5kr6tg8Ud8VjKUygZWjk7I9KW6/uvm/cdfU
ME4nT99jVmRs8Lt8PAhoOgAs54LJGIbkTDXyFwnnbQsI0Ac085Ma4GhccE5aMHSirbTidb1WW/Nx
09cVrd6ubiTLZCjcMxdaVz/0hF+nzjTptQltqlmnNi8dFCEobm9T0L7ihHyCzVc/WFo8XORfeSfN
5rorYtwKPUtvxk+DkkaAkNeV0xC0xQfmlvtep+GaVB/m1E97O0fcWp+S7/Ta/ogB1jHnjoRQvHNQ
0DqqSOs4CosOAjHtH/3Mdf/iMB3kJS+VZPxpHxLbHB8SvtO1dqWFs69szbyNQApdxiij6uK7u+Fe
fFUzujSVJHJE9EczPJd9twJ1GWtJSkPEnOsX1X4wfK/Ebvrd/ekc3azwpfsKfV0g6/tuaPQzgdap
dQJUjW4ZsZs9OVhLfL2tQKYwNoPM/s+ml+3v55N9b8E0oWNOVgqqT0chLqUA4ugrJ9CNVtsOhi+N
qwYM4UqtXMPJqJH6A49sDu+mk0E89NY5PU3/koxXBS2w8lfUtZyzj0rv2De1N4v0jTuw27e0+duy
rq+50jrzu1GZX1HcM4v3JFXmGkLXVqNgnHwzfVPrtdG06IEpgA61cqma7eJXIX0/ASBCPBCI2OFL
MDgkmAAt1vZ5lHxQskrH2EbHd3iVeoiOQj24zoloEPKQBJUxVs7V2STUNabpKvmrxDVy6qdZyC9C
513V7q/x0/wwAv2F0YUc4INI2rZ+V4SVYvft1sOWT4+rBk11WDXKI9BPZxw0thi4pN/4Y0s6rN+m
3cNFcm2mzJ1R6S9NyhETgOcZjRTSOGlsE9N+CM16vdYeaC6whaJ7eERGrk/rPC8lG2lmVmQ+hh+u
cYzNw2W/qV465e3dctCxS7MDv0ScHA0JaF5Irru9eWwOSYFZcj2y6tDREQvG35DUO18cppyHhJ7K
mVV02aWTHP7graccKuedQCWlP9hl3vFwSGDxWCkW5gCwq6o45eoTpVg9IoXshgYtQO65yBrLfGYV
Dhs1idIe9ZmLV8Pl/qUMorRWFnESkGon4QkVg857PDkevsPHfspzpVImJ2SW3S0k3ZWBhzbgQ3Hh
TpDC2SwsLDXlgpKPMuekyZei+tuaOWu1vituKqWB7Wv4QiGQtc4+qeSAtXAmCRMSNc0QJs92tuls
RQbIC70Jwh8Mp/lGcUUxrmVBuvLrnQKXaM7WyCjydRKURn5QVrwgvFeut+N8P5a1y4NtOV44V48G
aP++5+Dv+nuOFtL6su2X9T05mX1/FEtGxZE5Kc5vOXXLrJ0y2wwasvkXI7vn43nrj0i5w5d/Fmaa
m6uihT36079bAnBfRpqVnmz15rUpn92elu47vAThp2Z9wRqsqF5aDP30JUGexgp8O1eEa8lPZI2u
3bw6auxPCQfeEMe5rSdBaQ7yT9XwFHk4g4h+LrO+HCcr55iNZOqWm40Zw0eigPAeNTju0lxE0m/o
spKVtLds1guX8Zvt+LwMKtSqAxO3WXtNggC7IGfdDobIiBg+hoW0gZXzwWa0xtmKGH/T+7TAaK1T
GutDUScKpaZqaef6jEAazLI6ritCyUQQRgi3oUwPZXh0RXQ25zRJDdTTfEprvvhUlQjGI0wthiG2
/sUUBtZ7QAguRhTYndJhz8A5WydR5Sg1MNrDFUFvpM1uSFMPpbGQ9l3EsuXG1agfAaw5hdx6/ouq
rvLLlJuCYu5Qq0+Bx93LDv44pdkBkCsDGJzlxfkJgs46aKtYAjJmd97fTcrUvofhW/0i9NXsRKxF
9F+p02EQqMurHWU58vH98g7Qt2MzOEq/HAlBL/rR5/PAyxRqV2fU1ac3fVV8eZIfojDqNXJQtGP3
o7ZvkAcnxBGj6GTqOeUitBkas+hUW3Z2KHG0Q6QKYVZdhxklprpPV3QyG4ZhGYgikLidpz+cj7yG
OzV/d/4NA9sTbhhSssN8gmkpGhVIscg9psy+FX/2rDFiLb1TRHRee2vE/fCHeKB/6T2nvcM+JtNu
SVTOHJjrP2mEtHrvS8/oXEBT5dF1CWh9E0uZF1UPfJbyX0HHVzUROGRLsrQfBBdqHWZdtDnPm5oR
WetrDYUF7lBBmIAMm7b0MUg7QUO9DTaPBXq62ip7BqJUsWfV5KJKOFT+widPnBstDbjuO/u7Zth5
NZhb05R6Jt6B7p+gQWfBA1YNW4NLCwD/auaF8DkhPT0jt3cZHIQO9qi6cKKScWxwSUKxu8hKlanV
UZ5MymPVIIXzLQG6Serj+x2po4EPmZytBpF5vfSkTME2U67SoLkPhZyW2HzxgsyDBcXq2wepcSP4
Irkr0dcW6QxpL8EtOfgQbVaJezViG+P6qIgjObkqJ8DSce5PQ13xFiq0RGb9CrvwD8agGNrUShl4
EBOS2MEopk1tEqaPJBf5yZD/HwG3epy+W5FJXxJAvHgtmQ9rDP/0bp+KoudK1f9Bdfz0WB029M//
nfx1H3Hc7uCqEbWwabRiPaUX4E0mtg85zoNzlFfI5Tu49q8i6GKQhU6Rjr6EPJbLdvqjmBVlUfFk
Axi6Ivyl4TYZ3LygixAMenPJ8U5MtVihGh4Y7DpqkcDamKMblz+yUaOO/PKTax7/E+Z5MlVzzTRJ
1HVlca3QTWkenMFONuO/Ig6DB+ZBTKmYm6//wv6xoNIJKDQgJTBbT1PP2gr6yrhcTV1VOP9fboKz
FW5HY35n4TJVbtmkLCQv+PfXLqTMB6+zSSSWPxVClp87aP71j6RePq3qU/OBTZg0x4vmcTjcsvF4
iuVezKRmV2RHAJmOzTxym0xW190ZRQTLgRZe72zLQB7UioNB/bjBXZNU1Z8HL8H3gXiAJROPkK3E
872nns1SnoVAgZGkkml4C9ixaA7C9ji1iB5SbgHpglqNsIONyU9zBYrv/+YNZrtS24LHiR3kD7S3
MAs68fq1Z4oB5A8KZ+A2djHxFmnuIvZC3eZNgm0AnO69UdyDRaCbuzKkDncwPCGkmR+QN8CNmqdS
KOMEp7CmRKXnzdGkbdATm5v8zhDEYJlAxFyQiG2Nlgtev8JCiISZrR6DP+SXOp6eyfBmGalhWRNS
rRSO5DEh88biFSieY+mkDynnzLqnSrCLiJ6+c+BCj3H4RBgF4Q2qhSjY/qiG9NfyL6QRr+g+yDQe
o4msz3CncJo4IhGbFTdQNmIPvo9d7zH3yU/ios7+Ceq9zHKgxVrCLT1ChkpzDyagGbHkkySYqqA3
9WROzn4dYwuFG90FMsmeVeBDx6v5QePY8yTriCyJ1AMTgWuZ72oDUt9mvQAAP2HHbika5v9rwhf8
+W5ESHo8ABKvtoAiGNVrKLCKWb1onCwI1ceyiRwEoB/pu2N5Y9uylMlJktVRXMAK+guGLYlsVZEn
tIdbU3JRQKzNsZocJlk+IFYfweylDqUgpqzK7vClNj04ukwwugISN6PBAkchwk/07MGK/6BwQ+tW
6mzosVeenzjrDYtYt03TkVmGZCl5TCl1h+gh2ULqt6h1PrSJCn0ZfBJps9TiupK9ROrhe/6AI8OH
etra0PlSKdmJnQdtNYmvQBeC88Y0EoJ1Fkhqsqjb75WmCq2OUI2aiFA70qm198Ft9Dpkk692t+67
D3A1SAgxD9AJn5Kr03Ts8GXkh4LORtnU2xL8YdszTcI50AU3r3mSsfGsAYq+QRBXBgZXxkaSCizB
nIOgCXw/h2EvNQYMbVszJ/dvJa0A4ANeD+w2rqw63rOFGRJ/Gn7aO1PtpW+1zwo5pY9tTmwNgLsZ
7Wb3YkzG5+zgzxkdpofOl12Zi9m8MFby8Z/PSaeO0L/mvRzMPSXzuVvvBNBRkKYdOBEZBE6hQ4GQ
yi9vua/c3K+5EV02eEmEEDzYrCqX15mVi41P6C2fIwC13PJZ/8TIgV0OGYWarXyjio6ZeJMwxgOT
Fmbxv0RPkmqo6i4Y8+TGwDi4g+ZmtlHodye+TZY8zUsVmbsfpPCz1/dy+iCPNONtpOdXtkjH2adB
JT4htADBk/tfHHZClLUTEEW9tbhAwD7BAR9KSss3oO0KjeHt5AYCKG2cTgW2Njk+KcV1ViSqJcHB
/p6fzZ3sMSHyk1QTRJEjvT0nmdF87rTFYOncg383izEcB7Tdyo4Tr0+Br3nLT24chtmWdJDaWOni
Q5XFWk98VOzrPRU7pkcBBpUbffHnKYfBNG2sZb8a2ApEWk/4bdvwHE4EBDoggvFlH5lgCXyje22d
GIFp0pDxj7Y4TAsPfyY+4/R2ry7mA5pf6KmY7yKxkgneaBfLmO+8y+1k1UGe5fSViPSGMoK5pTFM
TcFzSLTW6Boligasm8M1YURKFKEywvqeRZvWPiON74sioorQO0sFa5CvrWsM9ncpzSpIAHPPWMtZ
MySU1/DHvb0Bv4CTlIxH9GtgDMJp6sfDaOQKKiSzCZp///WRofyQcS9vlk+1lvNtrmnvpN2LtXrY
da1/9lwI8uZRaSprE97YoB+vaioWdJR61hciZjJX0g3AujyVr0FBfJIw2ZBQfWiBP4TJPCwMiyjP
48ZgOAh4qL137f6GS2b5dzrmiqdBeGN9WYP0pEAhPiTxd8DYFK3kYMjz8cUkdhPbXrBRd8DRPRPM
Bux41Iq9UUex0V/WP3QUwKSarGZAu+LHT9sjL1PHjun+iOIk1Pl/GvlD1Yrck0Bkc2lpIO9R/M9p
M6gD9Wxnu0Hu6/E/mrSLBaIvTQN+Ls/8pY0BW9nGzDYqSzI0ylEEY87Chy6mx72OC+fcQcOhi3bo
iDjgMsSeTd9wZRl4DGCVRDqod084t37NRUprjTXaOncVKUhf4fllOsfDLmsB7fokfYXZvoUy7sNI
rK2SDh6QWTKvgXE42qN0FLmS/1twwR5/2+mDcT9gsKCFAWxlmib5QABCDHZrQq/8NIkLPAloMqE9
svhDHV2ETXmQjB6o910ZTDWolIOzyxP8CVf11G123jFjA6z9prTUAcYedIyAO85YKfWjwO79zMIf
3Cet/nb/haNvTWAqHolbMnflYYENJXOeq4zT25fo16S3lIzDqSuuer6Cpnr5lJwwM0Ggsw9s8Kki
g6BoecAa/VdQsClqka0bIcpgai1M3hogbbg/9996qeNUqJts/3m7ImJBv75JojbvgrVQyVYBjzOu
Xowow9TUBbqcIyCUBKY86fAg/WCUi2kX0CurzIu1zABIitSL9X/uRzHLUhj2d//S5nQQHFf0vLT7
H4862TeOW4a5pu1IYRVRqz59yCUwbmeT5ACi6dP+PQOzNTI1fH3C8DQklDSYDjVhm7zViBNECJnI
YXovkD/ERsKy8UDca0iP/EhiMFQd3ynt2EgBbc5yYukauJNQUz4TlKyNa7bQVXriv8Y4xuRsipz6
lO5yw7mPhZdqamUkliDHpFHzuXUxeLlo6sUJ956+T787eK6uVuOMMSVDTX2b88Hh1qRilfholkxY
zKRcDgNahN6TWPwnQ869CwSM4aETAA/eyBMMV+T68aRrXM79fYqJeb6ZeImvv9Q0cO28Lde6Mmgt
KPVGiHZToTNW4tUxEM+nXoxNRfygmgvsyL2uacStD7jPK3D2aiaLfPLZmOOgcWp67zrtZYOREEpR
lBKnR5eF0b3HLYtlOnAP4oSrnp/aDPFb/iii5pdtzsxeYBCl7pCO7s8Ze1mqIvlkKolwUpaUt3wH
FWwUGTGzgoZDC4kuN07dfP0rMwTyAqYziRFKTUnaERXmXKyvAreKVIk4mY+UvQD6Iuj+1n9TOFwS
jPlpOPy+CprQo/Wrstd9KhBfbdZgVhiFsqcpwEH43fPXT6XFD3lbV2pt99d1a4tTjGKQJA1eqtGw
5BtN1v3D7B11IstwII39QVreqpU/NwLuKr9viQ8nww1x8xGzj4Tizk3yaVYDAS64Cdb35fjKs/Xi
aXS3py6ucCvy1Bs/4SAdwj0hJ5Zolqzh6GwU2gX+inLhgeDXxKO/0wnDwwsYdopgNo0rIr717aVa
c0URUhZzrRJiVpk+tfWrAs4aeuLB/Uri626JqFNvru4Uel5qsSBN+yMRA5UVtBTWdBefutuAAp5o
Tcz0wpcQ3foXpgL+sfBBV6GcCLdyI6MENfh9HFhhGjfEWauUc2D+fUpX6k0jYcMp3bnPkbkhXzPW
23gWlwgmRSeM6k7xud8nibYiWyG8moCl91CvNaRztV/1aT7gOx3zk5D40k/jlj0OIy6SFkM+41T2
fFw3RCpPtNSh4PuQke1QTFXn/3/DeHHmy1AXHlS+Z8rKmDpoDT9nLW6fnW+39m+ZWYkpgZB61/cA
V+Z6p+mxQAhHrFQdmeJwLD+OJqLTuho3jKD5Wy83e0pgfIPuT9QMWg8nNwKzQc4yndnfTjWwi619
380vRLi9I4W+9G3nGSQ37ce572M2KViOP10VSn47LJ+R7Gb0LUc6dF2Cz4PaoPKXgLX9ZU8c15NE
ozHC2o3QQlDkfwgzh3VtBBypGHefrLoNZrDsCyTAls9AyklRnL8uu/GRXG470TNAVmUCgS56JHS+
Tg8ED/3XWpr8AZBNgdZnxH5K/Vmy/p/fCbCb8tv5UXiZJCkZ6TepOkFrqKqmOcep2HH38Gezixk3
HH1TaskJ0YBumqoAr2fxnQZVO03/dYAmOqHlM6Fyp4A8l74RlLF8At8xfruoevysTQbQXSsagZAW
wi5QS8LxXCF6vFQZfmbKK8C/kvgzftSpI1rv6z+AQQvuH+dJbEhbhZApoFxMDzrc+atUgrrhQNiH
/Uwt9YuOgT5oTA8yQJFmGX0yZFa1EEK4J/Tli31uis77e+NG3yDgdU/tWr/HVzHEHw7JM5ryqAJv
p3yepZG8fN4e9tyVkqHCe2q72M2idknDyXOfLLuc1kJnTyFuBumPXMbVPda6HYD+kmQe+VJRJmxg
WOquRdjDHrkm61bq9Dp8CCXr5ytrYqfmPmjhyWmn4gzs9HVhZ6qCXTHzPkxHkrBdD0wCm+T1bvg2
e25a3OX2IipR0cffgOIoaSSTYIW05vEeW3l3K8deNTaFqWAt7/9s+nqJ+ITCkduSPJmhDCjf/o/a
JUne5tOUZ8cy7sXmZUUpdwzVPDXtDwM4WxTRKuezref35/70wObn0zRxzGsHczvByJOkiIp/9Nxv
+mNBwdGvOcNhb7lsm66bpGp+NjJT34K5LtRY9QsdDWvVGjzaSDy8NOiNa6GztAKDN7yJEfizCIY9
U3kLybinrQBhzQPGKv0jdzEGDc7Z2kYDvIx+ZSrgsk4J70KGUEb1KJyDsr+ewZc3e/10xtGOk0O+
e4dDs9J8owsDBIgW9pcI9zZ5W+hq1Rq31pt5HVb9eKBjW+Zf3WCT4SDm3bzDSYV9s7rC838kkh26
wUwHmoxMc9vlbHxaYJBSE5Ntj2ve7Qc4PcbDQPPqYta0VItIfshKtu04G7bJMWexWiNOxqIlLudY
tN4uAQ6rtxs7g+ubCdiecJ4beSin2/6Mr3a6Qu+yXE5rJba/wanqPJYLjZy1HnscTQ+MJ7DRdpp/
EpwpexKzViSMraOou1D870spL6aL/9rOw+1HuVgNYrqhiNug7boCj79w36vAzutwI9b29IXqFAJz
YSYCMJxnkk8sgeQr9laPRKV9neHZTrg8TYqcKfSpvpLhO1WQMHMHkDplEhPDbTU9lRVNwsJOqZ8l
lY6mtPR3hmFiTeTnBdqyN1NqAeUzjidx3KEP7Jk3AZYalAb9iJEmsDogPCu7r5Z3qOV0Gb+Qt8+t
rueVO/ezv9a40DjbiC2A2to34Afloa/PXvzW0JCaouqlQIENVvKOPzHUKaftPZl7IiltGmaAPSjO
o8Url+xPgtNmccXIx2wRFhSNL48xjjN0NmueQ7CO82W6WD6IQ6jL18zs1CVgMfYH8tgQk+/9MSkI
TDaVFY/ecmAZQ7fb3P/qb/wbnqM7Q+zPOYn6sMtz74mds2P83rIwnOOn3jsNoan9JcJw3/y84qV9
oCNVfZ4Nbz7q1VLdNYUqNP3m87w5vWDp7mhpjdLlAyGGAgASpCg7IkTFFPyk/ZnNWavmgB/oVkw4
Osf/WyvtYWfodSPt4EvdOxGDMiFptXoecQVt1MD49DOU5l0wOIzNBiXPi3+vR5ReRTMPEly7S3rN
LnrcVsk+CFvnvx5y6iEuo1mf3EuwaKVXdh2KKRc+pkNlAW2HAEhUkQ1S+QcwtEOT6wAFLWWxN+Nt
IxkP6bAzZH9AscPU50+IALVJ3roG4DoQbAIzRFLpvQVx4HqSn8iANDiKBxPCWk8quiNPxrnUCesX
IouCXjdqrOjf7P69bR34roiDAVjaC8g+ubo03vjhAESRxLtfQHkiRUypIzdkRaquDGeWq/OB+XZd
OHPhYjWwCpiyfHMk5okCKy28BgzhMenI1P0vqDB7ylGuecTjWYSxyfOpIugcbA1/t8lgYu44RXxp
N0f6tQYdovSsgW9StQ9Lw6yTaro9naTrudX3htPhNVygC/aYH1io59/jTK/DxYCRH7YOkLYqsr/3
MwdqFwQi+3WVOMXPFO4G/lyXF3gl6xyiAbmJOLjH61+5bsLlP5RGIo0oZolECy4xoTnt7ZZ0dwDT
aCmUttFRuRUwwFHRgIA9Ch5X9OLqR+/L/gfWgqc9okVnN7/PTwpMJdY/fydNHmHuyFWrBIzm+0b0
EXiFYPv0xB5bPqod/4VY1wnihmQAv7enAs7wDNYa1Me7n9pMkOHP5E6t4vSWMsXOH24pCisP3b3O
UgVBa3B4wrWdd+0zkZZF6YY4fFxjaSGQ+6xkmu/UAqsbnbvBMRRN1AoWeGH/dnwM8NiIvrMVjPht
Fw7ASRbv4wg+NeJPyU9mMM/BmmCWMRrtkJMpZoOvmlnwB/WjXsbptOzpjnUGvBNnkvngYvWddbTo
rgth0GjAS7J+A5trnYQRRgB0QRxNLLTyNPT7+VJa8PuXaOwFNjxZXaEYJMjfG1lQmFDFZdy2V0uu
kkrp1Dd4qFYEVvwjt9joKb7rcElhdUM9N1M5v5dXIut4xJsgQ7lpQz26b/dWVeiuciIasHzyTthU
1A7ZUO4NZdz/U5zdZPqWxAyhr1d4QvtIkE3iF8w4B/8eVVYHLDn1K4r4aoQ9dIVDLfmrdnra0XOM
wnWgrm89HTPxYWKx+XN6BW5oKuUfYC2xx2Mgzw6gl7JR59nJPibFjfkI4tCdVTv7PZAjGBlx8snY
PcqVFkOCa6xwFBZRjMxTJCj5GBJShFd6+L53gLJ8NbVNQwpU0uNZKrE6ODIvVkqnxZOl5biOGPXz
Ua/UXLsUwgNH81d+EUWZr8hHBPck2cjosUEWPmIPo7BXUpGFReiRWAFp8sh55cb6Qb/VnOzwa6fj
S+xYxImunRnZlNaftBYdH9UE21tffT0zkT0MLtbeIPLOghajj01qdZrznAg2yPECbDec/LUt9jBy
zvAIxzgLqpg4uEnyuJYtEEGt/2gg4ZANPGcSPMVpywaY63I+9hNg1Cf1nUqVKUyt4/Vf0+jKkuoH
RB2FhXTyhC3ND2JbgLhOr2l6TXdpjS+h4MtjpcAQvRo515jWIbz/YfwYYPez/tdSMAwNNJdUFK0+
arbeJq8MznnQcIrtrr7BcbqAYRi7upxyRZhpWujaYiuruXxRiuHxqRgjCYh88KHi1xtQVR4JiUcz
1FDyasuanATqmjNy5wSn4ymqSquirxfurBP7FR5AMfLnhfNUrNgYA0b8dpNe8h5MWAOLNJVl9/8w
ZPX55PNU07jRb1ECbhsGG5T/hfgCfYV3bLeKSgDLuEySiJDxSmPisaxnjGHDnA7aitehiicdZQP5
MVwSNBKBMzyJixoJzWtgRGMlbf8h6ggkF+0+JIv89tUMpJvQSTTemF+96WqUAIbqt7xkcICpRca6
vZPKoGoWy6ztTegBQHPsHDM46LTwO9zonUzoM7znOdt4W0JSbpZEbQ86kVPLil/PyOYi3sbnD2U5
/Mr1q5+x6hhBVv/IfccOdthRVsvzWS97VpjIvwbrXHHy1GNrFnrP2HLSdOPdemGqAlU9BxBDxk86
kkAbbd22Bc7cJODT7jtDpIGEQkI1DoDgG3xme6/OEIyf3uYomcpHWanyU74wH2kERZiII2xj56yX
eJFTVIl2Krij69pyi/5oKSuGrfelaVQ/VkjtjzF/KhbezEk0x9QF5/shJ170PF5M9CjSP6wLDtPG
YMO2YxRV+KdGyzPBxtUssGb3WgJilXipviGlLI9/OOKvz6wp5O/5DrAbHpD2S3EHMtFgHKIEBlld
X0r4ujVRdhhBT6iujfZqZ4gqoaqu8seZeL3Xnm6SCo8NLY/D+T/ZX08ugwBxlJIdV7gon+RAcITr
ovOIpPiOpImq8mxS6tU+rol2otlGMxwL8XtAwqzuhJ333893GBnExrasD//0Qux+8V2jmRiXu/CV
YlouLGkjJOPS2LoLW3TyT6HcyMbJIDJPBwjWsM7lf/OtiwBxmJfXd5Lhsn67OAscUTOhD6PyhCYP
jtZ0bY8A9adVj/LbppXygFMD/wlibfjsmQRCFd7/hlNJcY0mJrw5pcVdp1LJml8HthIi5tw+bgFw
R4986RXhB7p+6B3YcljSQaAhAvYVCkAz38fnBI0lubA1rB8HrR3VN3s0O5oRi/Ntzi+uhbx+WEWr
m6jczJQpf4u5OL5tjI11KfNMNHoI8LojpcyR/5iOpqLO1tUvI29HHTdvQb/+UnYG9YkgU9moDtSo
ktXqmM1XVpF2F0YMqjyB2wUMxeCtvUPfmMc6MDmNAXRzKKL0oJY3xx1f8suZ/P2W9z7Vsu7+Kg8I
EPK0jdlxkh93U1UZ2NA9jRCOpV3XHjXHnk6723JJ2JLLpsebLkyaq2bJYs+KrnYOLgb9yjCV6O1e
ghLqN1Oy3Gb9E0AKGqwsEvdVSEnxYnkYQk5JQy10xdPDF/3QzmrlCbiNMXFAk2nnA44nH/9kDXsU
TGem4PUQdYCU9dQDPobqrqLlHuwJVn7J9wvXPNRIl3CsYxl3q0ZTJ26IDcUF18jtPVJQOBc0NE+0
2eZgz1jtO8beIZlSPCtOQnD2XKpO5LTql3379N4DAr5WbdT6yVn2C3sn3bFqaVE8bI8wf8jWn5O0
yXXq2b8q2X1qXuVMRFXL5M+z8FPAsOwRVTWRN1H1TBBPcrunVcg0pU4hWpUyIzFqhOMbUEP9xViu
/vfM8rUxBwKtQgnEf24UzDOK01W0cAL62LyHMt5CgZhv0nkgS7syu7CPW6twM7KQh8kZ3P90DUki
089QgqFwXN1Qf3YfyEh2vS0yaw8qC4t1MIb4JoV0gCkvUDd+ulqCcToYBCx/opgD35Ngbt88bp7g
vK8ca8q980MeN68oKpaW8hfABDavhgz7J8YtvRzur5iVNCuMmBO/lbbNjop9hmDV3x4y9vegSwEX
XtDoHYErYhdyYIZLLT/uSu3rIkYLlqwxU0s/ZiEzUOQeS+NJ/yC9yMFtN+IHuGIeho2WqsVMadzg
Mue1Yv7pvoGKFXIisEonsO2LVjS9dVPLVgZEYp9meevmO7tZ3FYLpsPue9gBwaEQsH8FedZiGYd0
TpMLw9bmjBc+SWh6i9wmZAyutPkmozs5XxkHyuRam8iApKLhGfYe4SlZA8idwLNd6e/tVcqWWs3S
oqTrkI0oEb36K+p8qa+XcJCo2JecLRtgOj04IC3cW02ZMTc+hkPgJtaiN4OkGQFzkIjzPcghhCbk
eBkzmYUmjzncIz8qjMxe0TKUo8jts5FjTLqnnk3knJ9A2FDPUkY1c6X+ybje9W6Ut3QrGpjy9vQd
SkvOAtZD2dT59xhOx3KBUjPxNsq/PjtFZYjbPVkHfG5pvALnzzwYNevqe3o2flaUQOWHFXZbWZ9y
fWXdFCKnIjhSI/UZ1BzET5mZaeOXxn4l7kuGx17ticoN1qb1RbsXhyaK2wITE4bR90KTDqCsCPLw
HyKUNYzVn0cyYvFvObqd7CJJQcT8kOrFo/Lh0xYzxWtfmYwyqwJOhjpS+Eb25vIdUy0PRkxJr8qR
vWu2r4UxxecQH7pojLVkk1jpSYQFsP791trhCOrCkPpJtHgltUI0qySmuXKP6Pa2f1pqfIoGfzBr
VI68UnHOT5md++F5IfxrDvPhyEdwNRqTjPXCRtpD2SPDfoaaUG2mBW3yj+cN8/QSDztXAXS1HbFb
O8F0tTX42VCOnGzy0DiWDBERCtEQQCNmdJkJQZxT8axViAni58IofqelBI48ytVa1JFPLivS3jK1
BYY75rx/5NJw5SSkxtRK3GxwF0gK6Dc99yevonuCDCIp5fkJ1ul2GFSCWSvpj61uUU81v7TXSEb6
TUj2xcx+10SHKzm6KKzj/utKZTo4CMcROLuQkla5QDeV17hREszPSVh/5Q+H6KfOdxlnZNnKFMGe
DcQfz7bAp9j6v/BXbsJAD6s1g3OIkLwXuZ23VN4cnED1+3ZwKKZKAYwHt2BoZ+eAiwwUu7NH/01r
wUQ4a8Z9a5gRQZ0m83enMtu+JQykbLkNFLDeTmu1grNTeyDTXa03hFqE88txwc++ebWXtfqm2SOV
MErNXr7UuQXGCFTbgDZHt2gnCkUmgjO7AL4pAygE2f/LwOXg3Bgu1FVLby6kPK7OtCng03STlXZK
1amnNcVHoBIQV/FVumJlV3QAC3VNlHpC8YlY/L783PUMXA2XBHfzBZcVvGJNaB6EqLVuvxPJryow
aWzDjN69R0jDNoARAavNJZSyEFrNsv5qF8WeglbcB7Pp3a4ssSYKQBhxPzp/CivcrVb8dQyrSufW
Nv+MCOtmiGHRk03y68Qw/TiWc0Y/HHSyAjVFLgpurbovDaB8zUa8/pnj4a1mcyr1LGg7Rc68PksB
jR4XdEYdRz2UzpbyE58AHHcfrk+Weq2RPOD8k2wJIrA5HyazO2+GF7xpSAzPES6inwSU6bmI5axz
YCvPkrJpCnpTYj4mCB6c/esxW/HiCij/PjUEzNg0E/H18Ks2runEFtM+Z+ydNMgfLGEYdj3W2o5r
JzkYQMJpcE9u5qwvEfT4bfzGmOyJj6EtGkMBbEtBg7sdHTs1ansYHPEdrSFiU2radntcg87NbAYx
0kAhNym5hj3vg69SPMH1+BWsRhDqfJ+BFidaeQD+KmdLemntrpbw0KVpGBAQnYNTsHV3DhOq9hVY
LqfzWbUM/ObrFUFLzcf24+kwJduieA3raYTUIV4M6NweQZf9eHieMq60DwBsXn3NLLgPwfop3OkU
GXcYxeqrqCd9O1tV0KZCtE6+l7zUXdUcWn6a/MNj9HiwEYHRt8z3Oy4RK9PRFNpehKXD/TECD1HM
R6CBZsFY2HKH6Tdj40w+eAgt9qtUbD+o+mJxdS2paNfFnOKD4bhDU2b7tv59lBRZrnvLkuijsjBO
tnr6DiG+nLj49hBf8B4vA19JXYkNzL2q5jnAPWRlfvrn3QHhemwcgnwTBH95cZ4kYfS9bT4wIC/f
/n0ised9H8vAhYWGVO2g8Vhn+X3fd8GYllLyBsZQj8l/5d5Bz/M1wjTlVlXLQhazJ6W0XC45oJb1
mBOHrmU4L7MIAoqqmGmXPgASKbz7t96bH6lzOML6KEXArbHf3H2KhyY6D5B9vlBnTjkKkB3IFrlf
nuFfkPqx7Cp3ehLPIGj9xy3W0rVp3IQpd6ZElbgNDsoFLviiTzdm2Qscwt5xoekopgwvwZ/4NsEF
g3XOsDeDaSY+Z9qBQYHCrE9EcKySZKgovF+/3RBkV3f12OYd6vTYjg4LAnR40yTqATCoLAmiq4Mk
ZELXN6nNg1JLbciq16OgEAyQuT8NMaYK8iCUGhwQWm0C0TSsMMnT8EJCDIio5KvSKcmodjYxk0Yn
I70hWAJd2VZwgvvmXR8y9m2AcGFpTB1KwCvFG/2CP6Zc34CAa+bgbTnevncjQ+IphtBf2uTPflGQ
fREGKwL6nUH66F1HXqDkpxiF8bjZGa0CsTkMJBLpKbhTIbR78y0ZBlMy8w/RpgY+M4wqp+ErpKMQ
mBInNzpjTuL1TIAQU2KmlNDcbEbJsgTCzh5kKuVRe0GjO5l+eZppU+oZVi5jUx2k/bnT8wpKQo2t
sUklTVwNS+Qa1NklpTFeRwC8rli3BKuVyYU4xzi2nSov5NEDu5flWz2as29VzAimS/bFnMEiNIMc
1nO5VtMFGxOnb1BjNQRoz2X0qEv8qVYXD3uuiRar52ThiEBNw90JY2epeJUeGUSSMFQJrp1or3n/
xJ03Z3Uz8cF5keZYgoQ2kOiEmBHfia/YtV1QE3Lhz7FrdGFyJ2fY51a95onGuM65Yk1L5hhof19p
VsG5+bl/imQKpTYInxD40ENAVKGikHFRFFlfdzfGaMsE/2UU90siSKANlS2M3q2v0T6nM3fTBevG
rPhcDAUTVcSLANmc68CtvxIeT2eRzqfIhGYLnCtJfOJ0QEAKfoTwoHCSq/SsK4vET9elTCZd8pb5
MuuHala+Keki8ju5ue2bw1KBJnnQAUbWzwKQqnanU758QdOPzdkgutpLSsCwjtAAUe1b7GhJR2Nj
KIFvNf6pSPvP+jeAEVKU1fxGyl8dtH2S4Zdw26lzJeQmjNnhC+E25SnPI0cFhHRSJPg/Vq83JU3q
vJusHm7T4h0/YuTIj4Tbs2ksW139UNypz5eMVYFPplQT1GTN+G297Yu0eMR0rwuwetXGqqRqzqeg
LtF3L1A9DhDj8owMpNOiaCQ21qHcCkTl+FKFm/RjMXITVOUNM0Wsw4ETOpXLaQbmkU+D2BY6mHmi
PMlq2nd/AjtShqbOzjh6bmFCbl/1da5Xc01VvjU3QpDwW89ATh8muOXxzLcMjzIPP9M0zmPlQ8Hz
1+O3sJ2MmGf4k9dViu33Qw+z7J5vglw7Vh3S6X98RmACiaQVWZGh0qzzaZUWW8wAx6JBaQsTAlIP
p8Gb7zNYI+v98aPpOUoQY3BcKJahResNmkneZULKxGSTrKNUxzInN9DUTV/Dbc2s05aKnTlCQjii
cQfNB80U4GPZZTO0laa13dUjTGkOuLZl68tdjpv1gTg2r63yT/Fv9TZFrVzmtSo+Ckzcvj/AFVdY
5PliMiXMKOgJZ69Z5g1klzFbsUxCBneoZXoMxp9JKZ+3/IMo3+Dpo0H8gkwlbIn3JOSBO+WpIdBJ
E5bLKm6lNN/E3qEj11BDsv0wobN+46rRgXJVN1riEIiPqtFmztawT+HQ+Hb+D6OvIW1N2tAYDDRk
gNZ2Q5J3EHz/bXdaloI8LvUZu7YWs1IHDWqpZMWQYZezm4TbOaDXvMn707CI5XjxIx7EUSj6LwDg
McZ17NJszuVDTYWGLWdesGNeknup94sB41flPPoxnD/cvOO77TdRmwT82ThM4rT4JsmX1xqaSSeu
5N4okPb97yqzXcIY/h5VZ/qJJZJGeG/qrLviJunyT9H+WCITKGh65++KlX0mKqyf+Sz3qO9aQRaT
eMDCnsT8vPJiN5x4OYSEMYKNc3IKa7z3tMPatbielWSeL+U6lJ2MwYKze/mdg8jzJaOgl/5V64jp
vb7pBEkz3425FJA0RXdUdFtz8mf4giBp/A5ur6B3Uke9uq1dMBBku4ZZ9NiareNjD2TaFsNvFBPF
rhFNI4unKsH5YHn2SNRNlWJhMNaTUT3adRJrutvfYKJThQd7yVjSaY++JVvlaF5lfkrg2K9VvsFR
0KZSwQYWBDOFAofqRvPYYUceHPpVCgas2u4Ke1pLDxhS0GWtpEDaE/Yl6d8nMZF0guWvMt+jFeJR
6rEpLc7EaakyB/Lfnn/x3OoVUjc2gTTdlvdYr7pJ4+aZFoIM6t+S9dakuKfqKJkpo1ZfKwu6gKp9
gcQyCJ2AlgNsbWdPpqNdWk1gGynkdEX7kj1eAAJWUkOBO+ZB8LCncXRT6cDJf0MucadSDkZ3263B
8XvgvTROXrj5p+Rm2+oU3FEm3gG/34RkCxlX+XG1tjp1ZGKOL9N/c/aruGs7WNgSth8YNXpv1tPw
4GoBHqm4nuP2me2qrSV1DY+HXezo5BPPL0Oc7tRvQxxRIOo63xDdc72dyrseZpQ1j2IFldlDrgtb
cRV+rNXE9n9v5WTWAr9HuVHb1yLr8wY9YSJPtcdl46gXlw65zK4fYY6h/uzJy3DdDUoPTdDLtPVU
hNUmxYs1sQyND++P5ZbLToS2yyJYBLzV3PfNJkicot76Nw3asjMOXhcYr9e6RkS7KZL+GX0vjbUJ
fmAGJhkOBeHyZk4bPnx1yd2EWMiTeqWvpRQdUuUSX8QzR5yLEz+YWUe5Dm9pLU11hypVdZf4x+5T
xhJPXkmLWpDPCs41sjtiFn88dfJKdzlR6Oz/xyaTRzYVWQVaFF5Mv8F1o4cGeyPELVjo1OQ+dQmH
hQvKZwKGxjWbWziorfq2+MAwgNrjjW3/ngXzYu/BYycNj+5wqkhyD+caTsnWv66OkblsjUfdFTBL
pKdtmdtofwMQzSmQtfbdkw1XWwbKK3wtrsKMlSC4RbawDzEytabuBZr9OTA1jU3nL77PlE0G4Y2a
sjAfrODeUd5Jezl5pLaz5APWjAyVM44/2a3vZzOPNHuSzXtpj6MwzYNBL6fbf9oxnIY5GyS31VFH
Pf4AqgTP0TGqWnKyWCjQlzOgbSOmH6qimWaiB3T6YL3i76NeDhVvhQakO43/nFVg1Ajb6UiIbr5y
y0zD3dMEyXNXd8qAgXvfiLSYHZ2bnuEbRGs9qTmBKNDcamwsKNY1l7x87CNH0phYNJdeGFKMwNBC
FYrAyGI7K3xM1h3sm9umi1NP/CCA+cQ7pahIv+ndZxjtOQtn37wtcLcp7z8y/ziJKwMglNO3iEVE
CNrUCSJHlNQ1m6uJ9JJL8jutGCrKR1hh3chRvwkGx96/LJl8Vv9kBgYBDmT2Jix+BYYnQe/xqvB/
hLI4DqGltG0BN6dHvhivc6NNjSpnGPaGt9r9Ky9Kuwv81Lt9+EnxFaDP24WD6N5RFkYsjq/9UrHk
MkrUydwOGB6tbEllQSOz01PjmlUkoS/JLmqHvaKciTNlS9lZQyd+LTDuuTA7NulfCU90aCyCEvbB
agIDKtHrQ8ovqiWezlttY16ckIscjCsuizttlcjRo4T5Cxp+vRQdkOq2x4lRxjtpd+Mf1SWPXB2E
DsuDIJT4hcZJgqPTFP7LFfFNwxbNmbTtNDKmeBk73EmIQFKV7rDpIiwIhr+k1E5KVOgR/L5ImgJ9
nzQcPNScVsqk1tpxBr9L7eqC5DFT3vSV19lwUDLWxImuAM6ttriYp4rn6Qt9yT1LjK+xEno7RZP1
E2CjK9Cmdi5SWCns2jO2t7YGGT2tWaMGw4evF8YQ+hln+TyZd1VUQ2fue/cp5Z5CLQcogD0ociXz
2Mp2x4k4+uMLGGgQJPsHIIvF3LkvmBA3lBMr45S2i1ZfdHP3Nr+DbaQrYcHiBFyU6LJdIByPWyQK
vTjBSqhyGvWtSvYFWsEXX3B/aYyjCfa1DskQ0+fyChYdTAxdMoDP/SiXLHQ4ODzww6o+A1k4wbXR
O/HqZbCh16U7IycXbamDgA71Xn9Qp1DcpUoaheITUjUtpVxPVkcVuRkGZ384kBmmhmtuRFBAjeMd
IVCRKECiXTs3nSU91ZuC/gzq5DjcTQJJ6Yfp408NtSsjhNiXmRpkIgwG+czWmIoOg2uDl+65PA2O
n90oXalBIQflv2G06eVCwHM/6yDQswwA/2MJ3zxis/WPEuerl/eLbI3twi6ZsRbRMGNXpmtykxHv
bORZEijsKU0Hymk3nFWWeHGOY7ApLkqpIGCZizy7fJRoaCaKQzR5dksDo3KI4ZbUNVt3m3JsHANp
8lBbkXbVBbwxNp7Nyeie92Tdm944RV8eVt1vzxnZKjq7H6XUJpwLMt2MTpceZPG7SZaTO/IItERh
odN/V6JOtjkcf87dimcVFNCshI1lVoPMKNrfag5rEiYdHuYRQdFNZtnVsMapkWU4cZMK7n2726+7
BGLlEhDUfe4HkoDLVv8dAqhVSt5lhafcD41KBwXrUU9cxEWB+LxNHbLL63maDS0Y7Y/DWSPBowxs
LEY0fcqfu8IFLWO8u1cxfz/z+EgTLMd3Dl2Wg527PPuBAiwprKn19aLz1dfzQHEOcuo63xCf13jt
b6TDUxZvFd4QGFt94o1eORze8Rn/sCu9HZ65zIkjeXqxm4RWA8MkO1uL5kMmyK+PsIsDMnGoVFwB
XrmXYfMrh9nVlqfARi4MFpwXQTieE4PuRZAahRRNZPGqdHyVR7EqJZaghjUkjfg3zRzxl8FnQ3tS
sn8/sPLUyPtSVLinERdG1Y87y1tSxXmrWbc=
`protect end_protected
