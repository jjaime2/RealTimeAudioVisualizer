-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HmwvA3HeVah70ni5QhZ+cnSm6bYfalvx9TbW1Xv1LM1dO1+n+WpRmgJUK3t0/6TRHxCF0AOzqEAe
mJ27LwX/2rkdjJyo+GK4ufbydtIu2REBcbZk9sRAO896LBNhrfg/K+HPEAFBBGdwVGgUhrA8OpoM
4dr5WiO7Bl6t1fK6LQDRddbOai6Dx1adDvNuNHbYbx+eo9VHh7fffXAjgW3LPoFefoobM0lor8zJ
EyBCuFTNQkLyPYnFfQyAEauK1tsCdn4BBaws+mW9hzEAIuDwSibEOM6GJfoLFekhN/3/j4/OSlsf
buRotWftK5S1ulVYsdf+0oq3dxVOyaB7DZLv5w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5360)
`protect data_block
fvMOe0uixHtAOiNkuMGOf18TVnViK7JaTeSz32NYdGWp7LLx3Md83DjV46VL0Njto3xgDZ5R9EyX
RBmck+eDl7gcUcfORfzwqGW1qhf0TrY6aPiJk3fOdjuLaj8z2Hd8716QvJmgANRnQgrE5BiCWTTE
RYUlhHnNjkUBHoMCR3u7+zKYrstHOYtW7cOJ21kFqtpcBfbg2Ip/pL+Ni9xpc0k/P6XuRNW7qLsT
pIXWc/VZ5ejOxGEi+064YyEWcG3w9VP7/ucHIUeL6JLn8v9wezOLyDFFayQQkcQocyf3LtPRyiHd
4sfS57MxZqeduPvbnulUPG1bsYRbC/KOoLD/yfgJC5OyL5YuZHUGkajFFOq5HH5gd+P/zefJWziB
cihV0ubhuYRfDf7ycjbuA8ix48NwiCWs+v20FvT1ZpRvXA3uEV9rzNOqVYq03bQGwV3jSQLX94f8
lv39oo1R77I1776TFc8oBFF9zV/6i0/uhV78eg+q1ImYXIBj/gPLY1q/KTxdpVXejDwuGdrOhRf6
JUqej1AU6vDWDCvwHHi2VWhSLM0NXr8+nkGGlsC0QZCutV49OimjJX8ENweZCvQI2Iov3mK8kxA1
8qYnNZIPE5GBAAtrIojeO3GQHZugjAxgpjGRTUkdCLFiOV6kkvZC4Tsd7uL1o2QSdt0Wp2rRw1fN
97l/KtXKmcOW66e6DVvS2YAxvi/EUnHHM/CjpQ02rmNmN7oWWEhD4wJ57BK1YWve+DAww+Bk3/HJ
z8GFVtDCm9w4cvZE6klz08Kn44sHdVPzbrJXiNIQ7nfjpuLGMuYkuoZZVKUE1njQ317KWyrovo1X
BasoEaO0QPhxhzqUCvZzdiH7muPOhVZGLo09K1+/1aSmr8jdwG8r1sdR5TdpAM4aM3W/CwitwKW+
yfc4knQQya0r2+pG0RG9Sfxt4rVexAMjig2jdXRW9nXjnp1XwIC6vM1+NBuWIgNO5U6XPn3IYPbJ
m8CskM6lkdMmXIPL4f64Muj11cUWJzRj7jw6hdiLtLIMnMNK8YnyJnuQfJTLo1JMhuX0h9XYPnn6
e+wpDA0WG4MMpK4aMFWTQxbATokleMg0W5vaLiBRQdPbJiSa8lAhhfxjyCT1dJxVyoCsrONl9fWX
UmuZJ2dhvroEk/RryGL2yFtFoTrzXR0BVioufFfnSkYKnqr8JFcqo1QkKaBm6Atrm6JvRabqQx7S
AdNrfie8mXHPWULMzKcZIcwB+3nbsJLg/UGmozOE2fvlTDxKPojY7JffmVd1mlJRGh5v804p42sm
GzzJx5oIKBquF0MZ9pqzgiFu+aeCP4/f1mvhObP6dc4Bgzlf07S4wbl7lhci9ficpQiN57skOfI3
fG9+1lhJTNk7UhaFFJ7Q50tThWP66lGC1CFIHw05ED5/tvrghyy4wbHeJuKJlvjmCDR6g6nLIdM9
ZQKO5MsuBmIiT/UB/nSqNRqpcww4aMrxAQAbgGDI33jLIsizVqUNpeFGohU9vMgi+kmfpG3T6y5c
Hx9zlRh7Vji+9hSgIWNABmGZ93Y7hSA3YhEwDIP+hk79bolndVPysBn/xh98VdAGcisH1WEHRTEg
4BhjoYyzRjYrn9ac0HT13t49DozRTzO0bQOdwQlowX1bfhxS/5yR6XPqYVU6OIyNsPSAN30s65du
0LfA67pDXb6fnUSf6xDXf9hyflolGQUBCUKZUK9LfqfHWkvsBSDXvmINKfEWlG7a2neK25uQ6B5e
p81nMBRCBhk9/9WmgCcdUogF29wztnECfX+er+4xQkqNDZpAIipiUtw2S6Y8c/TnlqhTO8unFdFU
NIghXSutim8jetHAhOWwiksb7+4czoLsRJTBMdUcYtG6JCoMMs35U0Ohvs/nd4uDfNKo6qVY9NUa
s3neYZHZl5D4T2AUbRL9yEoX6SsTTCdRUed38CIwhZ+yWFxuEBJCVIn+ekSBF+BjbBYFQV6Q+aGJ
VZVDV5Qkzd+s01OeGWzgI8DruWwYwyAMviiu6vyW3H2Ic1B6M67GzZy1IZzSH0RoXL1XMdHek3kO
Qegu+Vse0JMYF766/NXBcgX0WPdtfwPrNvcBahsLgANtUxXUd9dHpNxF9VUAzoau9HXAbDzTD4ho
DqgBpyp5mzoWwmZ7N31bROlE8+aQ3IdJxYstWEshk4iZpdRO3StX95T6ikoMuA5J3F3GrwZlZvAo
LW5cSjES4Mtge8RiEiDeWw72dTFacwci+VPARtt4fbkuDxinTHi36gc7CiGg0qjFTdt+Ajd57ki9
6oPNfT48MC4z6BI31y53pMhnR18YAzQBfVe8efWlyKa5WtrU9bi4qscq0FgOJcZeM842JO0BQ47d
AtDMfPTAPimlEzSg5OhLIQzl0L8nnGotJPuC+201yAIBYdTt8cLFl4pOlDDXVPExTJaXiB6mBrO5
OzAC0vsDV6rZmTdBv4JVA97+wvROAHN636DbbYFiD/NEjz9aYr/j/47zsgaqD0EcmRQ7XwSSAIba
ts75TsXjqE8jfBnTaWvEyIPp2X5HzwUwfk/UxRWDbRNWb8PKl1l2/hWgt0CK9iPjPHuv2Lr1xQ4e
CqAZ9pUJx10FRzD2GIqx0F/hmd5a7Zi2Sa51OQZ0Y+UR/VP84bZPeGoSBzQ1nwIRQapSMfOlHXy9
sxh9yHaPYvaQ3w49CB2CT17/8OaMqiVeFtylF0xiUm8ieaAxQMBU9W7pJ6axBbA7qy/nOqKdICEl
EQ3Cp1G1bH+sREzQmk5fZ/MDPvvhkAVTtSKZMt35At2w9L3+fuLBls/gWF8qUXvbQVoiIn0HYivA
Ex7UYHxYVIDZX7zXOrcrtI951njv7xZJSg1cRHQM7zHQhlXE+5QkCmCjRtp7WoxZww7EriyPgoFp
LEooit5eQnxUepmk9W+z9n5/+Kue2abaSBZKEdfCWYCCv4q7XjJue3zWR5ExWb2KbcflH+t/oKo2
tBHuxjozUNiqaI8ERb1lWKokXFoWYypz7NkEoM88P8rcoc6tpv+cysmpWdbycENLJWtw+tXrY9r8
4n+MaAAfLd72FwjO/fRR5pt5LUcvwfXnHAmbbhp5sBVMr3TDcU/V452IzfY/RqdjeRFFD1sf6Kjo
77W/Zt/LI/NsMk4HQ4qOI4kHjZD7sLQMu0ruXiWjskaONcM99HlkZAA3ifltXElnaXt7q3n0Yjff
PLE0P0DPAWdaAk99s2oknaAYrcbq+OCwrQOM18+hnSlJi3QB1dy5D6bCt5V+Ew1TMsPrRXJRHCsE
opR2Iq3KOdK4W2oV3MiSVVa8uEFYlHubJv5Iks4NOlFvTZYUW4KoykpHQquGLRKQId9xoR+stnru
UNqqbNPNQDl5WjRX9w2plkNQP5XdLC0wOrSX9Qi2hnG/nDZyhBNh0rSRhhhfPxBWNkGd52h0BzHm
Tr8lDVysadFkTkphvGauwevwv1/YLsg669HjpxmpF2GhPDnDDEx10dEGYBXVHTqS6VTGmw9L1lVb
pKdO6dA3QkNaCYk6/WiVtLzP3TDETZ4UDIn0xZknkeRIKyg6D9ivPOedsR4NLEsIY0IcNbeer8Dz
k1KkfN1M+b12bk2lHRYKQVSWSGIjrgiCsfU5yMFhUiopwtrfbduwNRBMKCQCfLeYu/AHKJX3xbzJ
6k7KI/t9Z/9+I4m/IFRDXcEjaS160cWyVc+rH/7qWpjmQ0gDNXS8S2LF+NjGWGCgmzT/ZKj+5R8+
egA1HMobpvvkLOXUFmWLZJ4GDfTTe1aBJXgdprNO0jMNN3PSPSyAGLp9UOZEdJS5n4/FIxC8l07u
svipGH2Uyp5Z0knFl7pjxP3HCS+5gOVJC8pJtqMcoNh9xPKIdiNsVVzTsfSmOZHS9s9illY2fReG
FybTq+7eIjUr6H4PhOfX9NYdVicT/mQRnbVHOlvbB75yowkF5dhLhQdMjUrf2bIkO4p6naV9j1gm
A8z7zOf6v9IWe2lF3mIgQirHiC3OVTAN6UTgRNrSIUEIXDSvmQUANRaSvvC360E16cfaSels6XLy
NhPLw0LwazDuNrC02jYsvV5hh/bntVXM3CiHhK4piMOOf3MfGpY6xYUHhbHK8g5TKJAJ9a4tp20Q
VcQaJKNzjEXQgYmlVTPAWUAZJzlsAxUo5zLWZehbSNtqbZx47++7hDdrXEKEK/iQxIpSzh1ksOex
YHI/yfMp5in3Yfbx89kMLuHuBskeRoKf2j4qvsgtOgYynn5bon7xT/EfqCMqhnwwY8xKK9btW8qk
gGQIaF5XXKs+rrpc+xmrSBgHL+BvoONuRet9qFemB+0uOkJLZiH4tNOoN8Ejam5lvmj/CQmL3rMI
NqLPxYocp033IzGjLwffCvRVDh5Sg964wWTMt0MR+jvvD2X5ZHKTydFQeY/ecIBucIxTQ5YLjk7S
U1i1w7YDprDn7tkNDgx2OvHGJqGI5yRY4ju8lrVHfkPAwOUe2sdIOy0II9V9ZKYoLGY2RWKBWcNo
wbsdnkJ2Fag5EWullTJ0B88K+jvQkaXaLfXGdIUKCIY99gpMaSS4RR5pYsiEmSdpbZ7ZEzhcMZJG
/g3sOFW4UP4QAzD5fXVKsiBcMYOrlHwb6H73ggW/rDDj4yhs0dz9wcck1G/Tx1zKykCjuTHLHlPi
ZnwQ/LYozwtYnuvcwN1Ws2+AY8NXqPD15hbEVTiVD/wKU3cz4H+cDCU0FPnd5qH/kQUBGrQx1aJ7
W01Odco5M8oCGD5HqxHhjLIou5DyOT+o2EYB5G/h+LieX/J+Kil6ntV/sjzl1IYLBqOBl9UV66Ku
slGov5jys6BkdXADgEAKLRCWcoXyEgwNxinjZYH5m6Eefsicb9YuEpXkIHAfgHn3T4imXzexbOJI
67AmhAnJQGgzpgLChnU91DIdpBP5xOB8KeCkCsEAftoTuPMIvDZGpU9bkhrOTgUS2wylm7VoPIQV
bjpKNOMwfJiqngBJa7oi8i5s9v3gQ/DVPh7nKVUdlUr/GzalBwCo3uutP0j2+zgF/S6Q1YJhsIZe
H9nOzU3k5PE/8UL3CI/ec8r3k1xtUHR5oSY2Fg3NC91w9d1EzmSqcJHv9iw1dxofaKNvBzbBaOWN
CzwEn1ZEotuSXn+dvyu03cCKdP+V1Eu5Bc0TTrgZa6Us+yjCsfyM2HVM5kVjYlp9BP4kmN4uZc+p
YrPOYzRoR8v3w9QpvIQpbiTdw8oqEquRGdetW0AagHF+qta3UYZs2Z+mkCDEzF3/S7Q1vqUMBFRZ
Bb4JCdm2PseS9QnOUOXCs8Q1nwl9WnNpdTwXDcF8fOMlpmxYs+aLwp/S+jr1mrXy9WKVWgAxeGfI
6QspABah572QNpkScX6WCGL0KtOhPegEXc4igSTobXCR9gJBZJ+Kj3RtkkSQ+c/ptEje0Ly0ei7x
FggNJWm9hdnVNCxXSnl9aww/P4buDxVtXKVZmpuWKp+uMNzIE0clyrjp/qEtfuKIkS4t6A7t4Umr
LmkWhc+Cu56d5/vvYYnlpaXjS1vww3KnsyRKlHrcW0J2uvOm6J0PpES6pG+/0V3ZqvgGwdhdYhGB
0C6xP/g18SQNe/9F+Hfb1/Eyp4lPE5rkgNIwQkdUgpZPh/hC9v3lWwn02g/cqeE4ZqJ0dzokyIqf
wD7pH6DgpZTSl5pTzhR+6158PoTAJEcjUBZEHZyacuAras4IcuoPi7y6E4H9D/kXTYD0bKnKJufa
BMb9kzcvhc4yOr1hnFqCWzkHmWbkuyshNOnFc4ztHE8DDUWJ9mQehNGBVT6DrBG/dY23xWLBQss/
GZt0zcm5oozpUFwDCa/sOdg6XvmI2aGi4Ib3XuyAgHzgYjgBfHlib46fWmx+wgAXZ0ExKTCg0OYC
6FUE+ZNrsR37XNjTSvDpsyvIPEVGps4GqQ8HcyV0NVKiLOicxGGAx8WpzDsG97LXMonhRPubegac
YkmCcaJMzVomvd5JUSO6+jxkE5yc5WrVui6jrXH5ZAOegi4pxn/+4ZYFnHaUECUomBqQYZueUhpn
R8HOsa3+a+mB9MSAscJlwwlQ8B64eZ9mL6JZYSh/1sQbac0KkDkYGOppRdN9HnQp9dyCpYhClYn5
eqDRWVChR4VszHK0/zNCzVoZPYGzL0kD4KgIxMOvfXhF4JL/+WeKGTWzG2ptPj87d2MyN0AUYqyO
SmSqtPG5agb4G+Y6hqjA0mYGoWuwFEEqKFEf7v0tjimJv4ikW0Cn1xRYwrRrGlgvQ/1cUdCdaWDV
vNAS8ZZzH8VvCxGW8bEnA2MaYcb69cLGh2ndBCiF2BPmOqwnnF/m8RPRP1oFfZBmVpoASerSHb9T
KuwYRkQpOeSEq5V02VO1yCmxrCPg+qgj5J3S1LBDkJe0eLp/mxbgqPfYauEWyyveRCsExg4S0SpO
bUgrPG9K5UpJhv7Oq64pBHX7g9kuA8QOvaa7q0omj0640K3LvM55Hd4BhMsoek+1WWNp8y+J7tUD
epwwLOk3bU5NmqA2dUb5t8MKEqABMPdZMEaC7XTKsJ4v48e5E5Slqy/eKjSq9PR3O6z7kpB55NaY
qX7qgqFSFg5dmvr3SNfCl8Xejn0ln9gwv+1ExW1Xv7D78Fl/U6XJK4+6XXlXy0OaPdrsWi1VwG49
0H1Do8fTxZxMCeck05+00CErWY8s3WDFq0CmlZCLKyja010bgtu0OFWqua2GAmz5cIzPEKFkgRCA
SXdFiEJo7WMGrCfWIQV/zvpotBHae9U9IK1y9SIHv7087Sfia8Zk+py2Wrz6bbbGsEUg/Li8bRqn
gv2b4sIjmus4YVf4kZfZQnSdTdSMpPRTjywFCxAql6TeFWEOqQkR8SKBOiLzYpduWZXIoYPwVHBf
USHjOPtmQXYaLRPbkTJFA2VMS2IGsdCqrKDtWGFodbc7JHyPo8PmvhmXl1FFaolM8B1RkyllHSAU
QltQbULQvwNeBUkXAJqyCVuCom+oup2nsw9hTm73sXMn3V8FAflH6faU/DikLFSCmbCLySOwd//9
6qruXvvTfshxgBtUiC0xYl/4yjqXhFtNdTIbteiivZyoDhNrTA/zs4qLGgKV7FP+LNU/6eqp3ZXV
j9JPKj4b8gPVpxnFQhMtz3NOHY2epSeZjC2KFaQrS2qzUxLZOo2aWHVAeUILYpJX6zCnu5MM4Yid
TPM=
`protect end_protected
