-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xYeCgdgSIh+5ztrJAbXjbz6YJAtgdQW5xkhFX/cNjTc5507jj1vLOa+/fUXx/Ikk26X6TzBsehq2
4Yf/FAhZqzPDIOE1k/NAWo2aF5bXCK1j1ues+pnqVmV9TU2C7mfsDx/LzNFVzME67+03EvoknQdp
lY9ytCB+0c4UU8g06d9rbwJcIlK+U+FjLu82RWE1HbtimxBzaQL+WV/4/s7qVGlsaMUC5UYedDpN
4k3a0ea2O13DA9p3gnB2JYNcsxi5thOifVeksS6tc+Q7bNd0eiVhq9fU2ya+jonq1zUqIsh69cxA
7e5Myv/6nso8DRoO8vRg6QQ1u/RPnuNqppPwFQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6144)
`protect data_block
b5/NnaMBWul8/3ezKjt4JJGRq32vrrFiA3iYjAolMQGN09oNqfa7KmMQAXtalldRpAXCBOZ9Ym17
LLBtIySoM4gBccbgH+U+woUEjeO3vBM5oUoUJdt1SxxlHlDSGmqcry6OeU1p2F/DBAN5y2fc3DMt
lpgEstUbADnVlIcZQfRfiAPE4j3/GtR1HyOIDSFxmbHNnuyqWwZCmPx38angI0TXbwk8W1sbkNRn
OFygu0hFErCaThMQ+qxgnDfW6UB1wSu/UdH8gORzeZkkjUIpi0/9dTJI/9oryOHm++VXlDJDurF5
z+okwEw8uFhIDVm5NHbKkpJciouQd1znhLMHUmWMUkMj5vrF2tYv+LartscX/9XaV7WiALkpM6G8
B2Td0e+HWi9BDNiC/YbBSrGPJnHFhl5lCPK+RA7rWltuDlPao+O+sIY+Tm9a62LS8oCM6IPP353X
ZtVEH4WjKXc8zEPiB1D4leKeegDDcjSVtttzoHSplfaaDtEXSuGeJW/ol9iLun7fLx0YQ5YK0w5r
a5eQHK4tOtD/KdhZ/HHPsldrQmqrKiJqtwvKNZE5PzNQlMYojK06Q6U6BurNZbwUxlnhOCAGw72c
DX7dC/ZLCEHkMDdBz02vXNsocC7Zo/Qd7tnqIrVEq8x/D8tcN/POMUz3pd8vejmKkfqu76sFKdB9
GNIKY6wEMNX8XJaXieC5rk7RjiL8n+LspD2trByUzu8uX08TQ4V7xtUFnaZiOI0cZNkYIrp9C0G9
Poxa1TtSoWRBxjwpg+RMtTAgigXL/BM3r2AyCD76xsDiDZbDbdJa0BoNFuNO9o1ymDFaFFjdrgIK
qSpfLVSY7jCejnCwHcpxNre6Z/AxtdyMUG7S6etC/bwZgmjLNuay0rcS7azH/SqP9FxuuhOphtRF
lkoEAuhc+vlS/ys5xQfOIu8BBM5MUpy8ZIRrxRb6CptwbUxitnUVuG/m+kISwHghPhgajLFR10bF
Q0iILeQFLDE79CkRB9yuMxZJR5bl2Z/Lxg31eZW8TEYBGRDOQ1/vzwG1g95GlAZ+sVqvQaOSHzUz
54WcUr3hbiY51nl/pN6DESguzcVN4ZEXfl3sVelfbziGvBgtzLcDzJJ7VrCU+g06E5FOpJBt5I/c
OKxRtnbo8E8uB67gi73sGfYLU3wR3f6BD9UnPd67QjXQyRmgDJM7T84FKJ3zdWqFp9A8Mguf+fdn
7hp+mgYyuzaTzLbSYNPd/Q8Dzn1/v1kMyXlu93ERi9RpN7eEzR2PY65+WEdd33p7ASA/JkrwpzOh
jLvGpwY8gmbNJ4FPKQCX/5XAT5tA+/Veb5swcz8/8djr2E/it16l6CNJkRUzAAlsKnFc6WtGvNIp
64WWuPd05ganbj/GPP8k1Bo0isHb0VKs7kCBiKJR/3wwGfkrge4JY5pBBa/+j8lKtvjvdZ60fuV+
QSVM9r9Yhg1YbgGxsXdj4n8FHyxfg/fD2KoceK0jyzVBasTEDf32nJZmbAIDB6J4OpS+wsFmbpK7
9waWDQykq2fBVRVNIpxDbe5JmRHof9iR5i4tLB/3m+MoFdMVER5mhlXBgQKzbgchscx5KvbUayY9
ogy0MQsQPyqt8gwQmrMSqsbuI9mQNbpb4izhJzzLCjn6OEpWkqplcaPWpCs9+Yy1cJr09NqIM1sg
pGPbEZQ4RR4ESmITwQ52Aqdz0V8Yfkrt/g3tvtxrb+dmIf70i3TeLduPYGu4e1kRXzhcRIcV75Iq
CGSttQk3pOx6zJSQTmWP3jnYZ3bUus13kQujyYpyYYMknnd3nnAKLAsxWCzbQZMNuTtS7MQBxf9d
HgGBJbF9LIRz6SCX4QE9kL/Z7HMs/rJHqA5pIljbRgASBX2DtqyleIcmiB6ZwE4hv9BjKKafXWKX
NZwFJyD9a2c+EE9Lw6z7NreJYdlh2LltE6f6+8cpZ3SsE8GuwlqOyeZdN3lRnonPA0hy8UsehBii
09oLUKKt8wuSneAUjlVccMovPonwrjhvei/lnSegbOkkoN19SuUQ75CJ3iwPvBnBX54IHjhilGOL
FJahJCsicLxBybsTm4vIwGxp2+wwmpRzGi+k28VUTzzWi/AmmGDMyygl5kSbbZiF/8AP3y5MxcV9
illU+fsy5STV5Q9ukLrLkihe6ootx3pYJGyFjCqxpvVapIkGtMasqGkahoqZMG3CavefzREvUKtT
9CHKYc3iwPLjiQX99bFKOelfdxWvFZ7o78EY1nd1rLMQtrWkcK5v7P4n2XcY5rvxMme8tKNyZvfL
sX8FCBQxwZFaMwdOiqx8GWLfJ4DncfkugwReHxtKZCB1fAv876bch/VxYHImFua4D/eH06yL5mph
dlOv3+ZfLpHGxUP3g48MbQUVv8sAnz5ThS/OdGaTKcB6xfViklDxLfm5u0/2KPpfRN4WDQwcUaSi
Ig2eBzW14CMvH1Gs0lejCcxh9Xvcjc8AXo7Sy4UpE7UOEh3VuaMdxzc5Ts5DzIQfvR5NDTAY3ue7
MWLZ6ptvFULUpEsqQXEFl/RtnWOUjG5Z2KqWC8EZ+L4O7N2vSmIpwiEo/2+oo0FFIZso0ahqcIej
UdTVhdvllA52TW64D4VPaTGdItrOTYDhf1A0MbWi36acAGFGbm4hfpVO3a8Qvo3PGZcacBBSo+It
tFAc9rvupf6IF+v4+IXpcydfN3q198rtqJQjjAa7TN9iRQam1sXLzF4KXRRzvDUn65GNtS/Tg35a
SKiN1ahIsAlsSGE3MIzfUVwSiGgBeKztBJT4qONBLwZ+Q7nK8zsLNZM1KdMkUUoHgwwIHfVIQjWN
EggJzcbun/IecGqAwfv/QqSJ/FlV6mCoDzngwxnmdda4KJjeztiepOldySo0nKpC1WaEprIL4SzY
ApxMzJA6ldQAmeGVow5yDHvs3bCaRdtkta3AlMyHBGcMH1i9YHp4QNFuVKrRXBV5a7gwM8QmfQeI
ZZAo4m0x7JBGNpHE/1FSezZJp0AJKiAoU+gprX5ilOWKkjXM5boQ7P8nxJPybNDJ1NTDhaGBOlU5
6QnA5MAIRVVJ1e7J9rFKkuH69O3qicMHMJhVlDoLhFpgo0iZ75pcB1EodxNx0Terdxo9j9AC2fV3
8nwoegHeRMbhkG6avS2ePzTQKKpbN+KT3bfR9p/yCyWtYnrOR0SqeaGBnowmeeTtG+6zI2ov3/ms
u2Q7ge8Y31MzB6LhQqCqn3jZ4evM5C08r+jCA++PDyxdGUGz1z6bt6TThvaMdaV6j5LDFEB3Im/A
rFFluQTzFc8UlakTDYgry905za2aBcuxGlW28qzyef19nLyjUrJrze5kIrH3km+8n1zRRm0ivjXY
E/5jIH5dkDzuPoKtCF7MdWNhc3eNc5hVBpG+DCS6iRgowGegbYLguCOJnxDvgBkywS4U0mNc/wRb
nu7xpVExo/ou2PIf5c1SwrGk0lrEbtAL8qNQGCZc/g9it5PqzH/eo7KJCmK4vKaa/JGStOWMP7h2
HYib1Y0zWQJ/96cUNh7Tu1WBPp59RumeVu15+UrN1cQfvikyWDVoh+LlEQpYLeskp/qU9l5Kbbjk
MpoX0ZbtaieaeeNn2svAxFKSyeYC6PkVx+sajA2gqizAcgrEmqOqdeW9f1U7SWPjS8i6Tpb+ls8I
/mRyqTQ+rzSDIwJqNRYKgyet8DmiUnxEN3d1xdaTd5EidOZgFI+ah5jhYUXK8ujfM1GULRusgLHY
IW+zEX4HchrQnNVmZp0KkJvl1AtFa8q1HNOBhuC8QTpDXeHbeXVRFkO5mAhLmhxlRTQQQEtgOsGe
mwXBTglLghX52562Lqb6LFCHZjQWDWiu5cnjV7ju9gL1SkwqssV2T2jJUrMY2tUhoZ9iVEsW5vi5
sUW2pvdr652T/Jt/Uu8TcYUSPN2BxNTa7pofNiC60bEKCwwuXVirL3qorMfUAU7GO1UiulIqR1Rl
35R0vqSPqjcgjZJiA6Czua1n+a3ifBEI48l6jkGO4KxsiRctWcvD6iy+wXsaAyKcCKC3XCkIu+e7
uB5qe5Zf73kG4S8vQ2iVBep0EUxRpcnSTgG2FcGacrKlmy4apmCIk1YaChj+YnLMsUQ5AafbidNl
/9oJW3uw/heiqmwpzrpCU1RskeP6fllTht0Ox4tw2b+0YwK3kgsvRtRvsi8cil0b0blrnmIoPI8e
NfBYi5P9NQYAaCVTqaFbB9VPZKyHkp/yZUdoPuKjRWY43W0qlA7AWiPjE/EkLSfAjF8FwpIVQ299
uET6xBHpyTvd+FGdcSUB1sTgXaYaE3RF/GurqEcDRYHquxjKDYdRrLAlwTlwxZmgjB338ItNyugy
zYtT9cXjVoOWxXLve9py9RKsPdtAUr66jcHSYSFAtFbuKP+UFwuIER21NxzX+sB8IQFAjZzzzc9t
j7NEvmujAK8BCIVefBxxeWluglSO5Q1x7cyFNsLc7DADuWlZ2ZGjFd+/67+MeQzpMZaZCROeRYwb
8KuNBpFRW2j6M9sYTl4Ip5jS0bPHxkjYV3VaHlvU4c8qfbKnHxTFYrGhXOcxJv67veFc7AHPclFE
cxlsLwVlQxj/1ANencAngOM51ksOFRc3i6RgaxFF0An56pIig/3hXVS5VQOWzNrpPtWar0vSLjCy
aafV0o8Z0w7ekk125PxPXbb9AgREzvZkVbyRchibmo/HcCKgqM7LJaO58hzzXX5xCvTrpYL6GlOO
BklFYUXkQ5sjvTif2A6hGQnFTb4X7zKmH1OmktglgKXosaeCDYTauq5KS3A1lVdfmA8FMbGAe+bC
lY4n8nW0XeRaKLP7lscCmjqIwHBDjyZbKIZlfTLGO+cb8unPTVfubhyYiRSaw4pskaOxgzjQMYLF
yUD5rtY47XE1WqYWmTDG4quaXfTd1m8aZdwzk7oytQR6wyFUrrqF+FVwjofIQASWydmeF0eW6OZq
FYrlj4sP9d4dU7XUDhefZ4ZBBrqPKrqIBmIG4CWAzHJE+9tCmmS5AoLhPkcvBo9ulf1cPKbY7nCR
P/WWrwGaSPTIuGp0BdUaavaHyC+slrtJ2iAfjV80bBEjZRKPKdacgmi73/VyAiQTd7QPCr3G6tMG
ol68lPCRpbkr5SyfsF0vljkqD/17Se5z4vD+OIwZOu8SP+8igFjxXbn/28oSy5CGpPhXNTcxzyqW
8g7O0qs/rKAEypoAgXMpfvxteqrR/4DcZsbFAqWLOiIX+M8zDqLEGHT0G5RL7ADx0g07CBXrupsc
bCxsaqOwglrtHLa+d4hMprBJBlQ57qVhTb/a3C71u9RZAId+4w0UVTPRig2Kd9sZCh+0jHrMEWdW
2rMg91kpPtZih3dfXMGswj8G9v9jcbV8pneUzRa0QAFwZ8b95AAwoglQeQX8jGhlkBhN5i3HUOB6
3XrFZP1c+uYfn7ZRxUUddaNRwZkifHTrilq/jbpNzgjkQOV+7YXXIF5P6Kb5Eyxlp9K/DHvOEcW2
NGQ2uHwHjxMRSdR+huU16d/x+qyDVnCcNsV1nwFHpqKdrMLPOylFR09OiyFFZkgtBhjz0w+bBVYf
Io9WlZzR430KOFtki90UZLZJmcUp4o+CEZTLvzMy6/gZIgqzYqDjku3rliQ7cJM/GJ3apVSS4GpB
Hqd1K5nJcwyXhkEiqNREhb/bevk7v3cgmOH2Q3kLQgOzVQ6IjTk/YZOf5GL5WxQsqxmtssfRQld6
5zF8PjorjiNPca9Y0vMSAEWnQiOhyojfrz2n/kVoT5/WUMHGpLQzyIGxuwaFNNuTHo54pG6vZMl6
LTqW7acDjBKKz8DppcFT/jbCM9R3cOAF1UhlttXMOI45IKjBPCHZSTveff2mwfCMdaWxaoJz984Q
ZSdD8+SbTuPiLKBRbEHr6H/HdPd1GsMQ0783BOiXCJHkjmn+F4b1t6B3xbziN7vLcRrvPeN5+HlX
blvRXQhpOmGNI4DcEI+ekZAfv9lo+DH9n1TzQB+Lo0AUO8uGYaKzNtygMlVrz2zBuBKzt9yDQZS8
CT1477XHDTpVk2vxpcpa/0yzx2EGaWQ4srWYL+aFESfOygLw4YopGdNDa0skbDIhxuQiusEeSORr
VWTe+rNueOKt0fPeJOWWXHi523hOVzx8HxG1mf9Qt+rIg/+Ilyj8FWos79lMfajE/AWEX/T5fINA
XWQoJOYGdzNpYaa4esxr3RBjwHRkn/mXutmc/2L7x6bYC5zMnTyeELeOSEj/PSut48RHVVqBzG6J
i0ycZIh+vY2Y7Y1EGa0hdrGthB9mjlA9uCUB/01jHDBATWm3upUopnA6N36EAgVAB65s3Ie+XTif
09NtERAgrkyD1nUQ1sfLwLOI5n8+/61VVWHHVTHevWrYcR4+spciIWhwszEVE/c6ObM+Sgvmu+77
oBBexm/0FiSJeE3jphcOaaleZYGYc1A9lEUNH3DEi5Vp2ywpeQkPvCL34XX7Iu4uterB+TQq2/r5
5LeffFMaFfDuV8vc8pk5jhOA6REStoX972E5wTt1sc4VXpaXaVp7x7LN5ALHi40d6LOvQ1Q73cFN
9NGfAWhjEwJPvtJ3l5lEN6e5ne5o1Nkmr9EL1DYwPaK9s8RhZTPPd54lEEwO/WqTIxwTkkLXOHrB
B8vqPrRixTrKs7ihPcdbpd0LjZVOR+Lattac5V7ltOTwukZwiuKvvOIck4sYlm8Q6vmLdUgZtChU
kIIAmItIvs7htGWOqoslFeEtALDFo/LKHPVU6Qs9wIw5pPY+G6NPIBjeUgYk+yDTGEW1xAA3HtoV
Lr97z75aBJflwiS38S3Pj76dmFZVrHM1dl7DuAVkLsSGLN+ekBMDgGFJXMV57sglabMTdh5IHMMq
djQLsqBmqRCzPJ/MNyMuw5vsO3jLTmVSxhS5UdnYRtfNNd09ryH2gP3p7KbSctMy7pagM8X/Bv3A
+KKZbwLO58eVXnDSFnvszKMHMTCDTBbVdXR1GjD68aePHUlLvZYg1cImp2a2IjpyIwmnSCn+KXyP
7EiTtj4p7p1gITP+Prp9Wx3c0qwy4+stZyNXjb2BgVb4crZuwkR8ryypLezwE/Bfpfh23Tivcpgb
IlAEbu1mjiqUDat3QkTVmt6T4bYsGkS8VsxXwR0n9gJfqp8aTwc3nEQJ11Szh5sx5w8lta6jEJEx
+6NAaVcHeaZHhfsB63S7ibZGQZhPjj+Hx8MqYJe2sVEDuuhk+cY1Q16gFVoUo9pwmbFKUDru7mNx
2MdasNc/lMSNl7lRdzoMekUZYdCc+KWJjtT4C4F5OfC+dCen3RJg3LZ40jda5YrBTEHfqYVAUMBW
nInPI0MdC6EKZy1/HYO0/wugdoFd7r5Ic4atmw7hVNLhW3JN2fyhk+V1LRgoW851nBHHMgAxPbRY
OyuWUHaPfOkTpZLp0SsM1AAquNxD3PNDhNEMaMd1C5wg+Oc+/yux2oQvVKPRgz+CMgxzFlh6uaes
IexMI9W4S0rZCvbUOCEO5XfFLd9Z4uc5LHMITqAefodI8+CQ1baK62iufMr3xz2T8Rg3oweX8oyc
NooqlHarMPei1Sw9r3BddZf8o1lqeim46WQxTnHIOW/6mMtlP9EyVhkosn3NdV5gIYN4nrYHEriU
xdabZL1ph9QAtZoinoEHndNh8GuqXMQ5Fyf7pV5U0MNaVGU8of2Ygtab+JaOC+h1m0Ni8jwx5Ku4
5xZ5bVusKalbTPAUmJTKGZ78mTJPpIVl1wPoSg2QzJWgxJY93GJeLA2FY+gbdn7LCNL/VijQ/1fa
LkgjqI0d/mqSmkEtJeqbXTJH/WPcXafxFwp4d9f4u8tAp9+94o4nnFd0bVHVbgCuHRzb3yEfOvcl
81tn9VQurwbYyXFWCabcbWANLoO6/LwuAvV7iNAH/Ps3OFZ7Uz/6af+vUHWHp14AzAAiYocIPs3y
c7FwSWQH0Ztw9qGKKYdU1CPrVZP/QKR+j01EmJoDy41kBoTf8UIU4KpAdMCNOS8mYUvDzt0EEHgD
hY5UYRR6T7hPcORy9Eum/vcc2uwL3pxXTMFJEvxoSlRiunq0lcv3Cd1bK5p3dzH3aw2PJDIQpMHH
swpjyHEHJNy3tpwyQwVUUvJhPZdpxqInqD4wOWI0Pd/QwpiKo2WYQZWdMFrE1PKcYov/rsTyaRpt
0nSF5VHhvkW8K/oDEXifApa6v69dah4ibs52ZkMbvvPn7vMAX56Z27FBJldV
`protect end_protected
