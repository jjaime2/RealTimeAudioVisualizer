-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
A18oGkUeWrCWGg+1tMNsxuLZmWY8K+Op1Y66y7M2B/HMDbc2O50pb/xbGMPtGmValLfT7L8k6K7C
EzElTckvsAh9Pv/ubXS3ziZ4mF9wPUjpuvxpCcD30ZwPp+4MWMabXOAku7gG2rjSzrtQfGiR/MQe
7VUMvcinPSbxASjLZFS6NvBy+5mFG8ulcN124HP57yo7BaAdwLINeLFp6mNWXURma9uf2KRLQ45J
WJQpyjnYrD0MVln1aH9BBrGodwNDh7/oabMGSAKHUNRQx0gr5fcH8ztLVlFxR6LP1Ym9lhNFJ1uM
y90JKPyGqUw4flRTSp2HIlG3sx3VOM/8FUDU/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23808)
`protect data_block
2ttOIrG4WTfrM+MVqPoYa8l/UJFd1sWU0cnkIu4V1r+mTcqhpcxRP7obRkKwLnwfhgZA0G2b+W78
RJMOVrbpvIopbn0QBbTw/sTYyuWTcsnWlhWauRT5BfZI0xqHXIOFQ6GjEaKTW898tkhiF4Y5XiUf
RXtktO52Ptg6liIynNgKpDhgc8QtElSIEZK9725kfRbhE3B31tfXFkPFLr+r/+zma2qGUmt9TIYP
sxIaqh8/MN8eO51DCQFr4JH95kP/VTOqgxIe54skupsk/dh9/STIebsdZ3tzw/W6iJq5G6FGwBjU
ywOtIHcpAR9yCGV5FfydXAGzvbRwz43VgAoIDzIMdahiGkioRlrSuiuVbuBi8GqtAu2tsgmmBkOd
p6AVG8+XkkbbNuZIyUzzPmnDqme4+MPXjXSpeCjb8a9CJSVpAwIIRyo8VoAt+2/QRB3vEgtb21Cv
5SyVBz8Vx3iXdCo4KhTIhLgEeBpFNdB7OY2ifMGFsmomJ4ONbeqFZY/vlr/G6u2aARUwYCVNbWez
gEzR0CC6rEczJ9LEYlYx+LYK32aYX8lID0YamoZhp7v9vdYkehAl7NqzV0ugkPuoUH9JNvl4yI5a
fb2K4Ei2hLOr2iKROMcdlx6M0qzIAkIbCRbLOgC+gwpt/fuTKBfMwFNxVzb4mpQeTtNAvZiVCSNj
k8jnclP2EpL5BRdJBzP339Kwfgb+WfFSBRVv745ah2YbujWsXMfPQGX1RMobtEL4LLxsCokuW5C5
Mj/2EQQjp0BuDSAtBvTqdQQxqhhpPt80ltSy09Y4+9y1eQCOGT3V6oMH6qEeI1q7/dC5/lsEZv8T
S6mzVhmt3ZIk7DxjFpUl1vNVQIzHaIL4ujgKsHOff3YSnjAmwl/Ev5DYkBG7r7XcTplydr5vVT69
rQ55Gj6MKrLVB05Px7qRWmpSe7IzndvyPSELPIpNGNpgr/7ogJkNDW3jOKUvHNG5wHzXw0rH3YYU
rLcKHDhTKvRVbBBR9//vayQpsj94QIwahWDx9I51iMYfHGhsz7vg7+Ghjt58lIhqpDmshDVuTdcl
2aGcDcsRW1ldvVp/UaC4bcI0oms0svDqt9snS+xkPrlkdAJg91KAOGG0dWHwpZBS7F8bU8feHPa0
P8ViaFv1sz5ldoAyGu1H3xaDE0L9vygpyp97C+/ylh9pkmDGLlLcdefn5vjhUUb3XYAiCW5EppYt
oOxaNOzUiHIslaSJvDLczDaG5pGiwj3ZIe3bMonaqCaw2fR05Zi+L7vHDLRJJvKjPzVe//LZ4aCC
2owiiZ0Mc4z7w041ojnsmYoaGJ013eqAkH9BwbvetqiXw0qsyeKxbARJjaHvHB3nz97ZiXlVxVFn
RxSM+aRPJ8/UWwVwP+qPDEFOCG56vtntD3boR1fkO6pPo8YYFjg5BlFITX8RtAE50dmUyjJIe4Tg
p7RwquYYLks04cwcx93gPkDsJSUEmKkPVZmlnnvTv2x+RQ+tISb/JKLzbJkHeT7CZ+NiThf31fiW
3LiGXp9AH9hQJIMGqRVSbwgNiRhyAq3+qPY1CUdY/gOnAFkXk9gimuNEaezZe9FeCQBHxMc2cnQi
e2MYNjKT9xEDIRUkP8D4d4+wA+84GPFoufpFhaM+aZxFzL9HbrEb35xPcdCXDA3V8X9WgKCmuqp4
IBld193IFZBR0FOLCep9UdYam4CqbqyADnC59t0PhgIcfIN38zDEkNtzIes9UkWr0DSEjiNOX3Bc
HkEwcLlQXkCOdkCK4p4rNipo/tyLON6/ylwyMLpoyVO+VkGn5DkDnFieGzg2d9mPi4wK6nEepTk7
A+66MveJEo+J1L5c+YY7kSSRMfY9DH5Kmiw0glX/P+OJGkLj+LPSbAv2QA3YKROdGzpDS85FZUpk
Qs8+CK8T3bkqqW9CPGExjfDNKuAuz3kQ14W9viyaiWViuYBkYVx2vDAjQuZ0NVQTXZjKtngLKiYF
pWQBAbnNGMdiUG6aqDgrmTlKvLmR9pskjb/K7pcesH3VFf1K4VS78gqEPgEbL3G570OpMhTNtzr8
vX/Nwd6gdhbWNhmJRgO7hz5qwz4JI0+JKM4fMf1SaF5HTW5l5N0kb8B4nHvOazLlyZ0DAaBKiLwP
MxqrFltBiWAlNOmDI9FQ9ARcJSgQuO9b3Y7qzyfAIEpfQGdwBQ9hDRhSCdhgc65lo49QlI0CPR+h
846+f7cgATbBiRN1taAO9vRH4Qa9EcprHQE9L7gCG+qqh60sjNX3a9JUm77ot4p5l9eErShWw/PM
QjJCz8NDkohy8u4S2+TO78s1q9+BA59Ry3x+HZuq97Nnaqm9kkaOmUvx2AbAkbVSgfcma2USU3U6
lYI6yf4xkDYNND85G8IHHAGECjM9vfdhbzhCpTGfuWw1rPRmP9dqw+5lDuNDn021kYLWtp/EYYJZ
Bjs3sWU6qUoHRsOChOZYS2tNQjcUVMPInuocsu4xPfGbsynTOy6CwVAreVxW2Sx/dpBkPhdAZNIR
FfTkzj5O/ZihZ9qtvKxxv563oVFN/U2JemsjQfLhoNB7L0qwFVzK0y74oqqWv3sefK+Pf7gJ7TS8
yZpS1a9fcfoy57UQ2nL7VSH56ayf/wmJqmgPOwCjlyFvcfo0DBPpFEBtmyI/mAoUUvjtvXn6Eoi2
UfYGUc0UPvuMV62Z8W64oSkNKb+fskL0mKNA/FxJzkT7R4AgNaWlbQvEcP/S86k+QnKSc8j6KRr4
y2bGIW/Y5524/xVPhOyYx4kxNj+eiExTZSfjY5/ZcSdBbwRYytPE9c3kUJgug22CoZX7RvkcRazK
uB2Ro4WqE6pT7Po6JW8J8zULpBwuJQU8MBmcvzUFv2kKxFf+H/AHzGzfH9773HX3xrzZuCDQ57HJ
/SMG3FMhiBheMdcWDjbKnSW/Gj+51l0Bk809B3hGzt6xJH/E07nndVaMXJgtck/Sfz9vIZ2qzkRe
Y7Td8xMLklJVkJlqTZP7Jk5sDVMRdIvDZnBj0zMfP9MaRFMCT27pCLuNNcORLK6cJg4rGbanxbC6
Hx10omP9C+U0WYd4JqzHzrmRYDSKAfXOxuFqGEyKKBKAHkVn2aEWvod+WSN3TSWIN7Av7qdtaAGU
RIG0pqiBqjGQEwQid8RwYouFirjaJtK7xM4WjLpwhp8llsbaV4WViVqf+ftPZoChVQaCyIf6GcZu
JLUAQzq5HQ9mRSLLTJfgwLT2htY4btzDeEP5LNxrceQJTXdwZPhD/CQ/OgbveJbmVoB5OK1spArm
9LkhmEt9VdsJehgkeayvmsryXBlMCIbKqvCEUQsOd+jz0zHaHr/FLEVmnzXaIXmgumXuFtQGtDOS
/Hxwgwc2IaUWUeGi5r1ldrSgYsrIbl+4I0+OgOXGpVSpAyY1X/lm5ywYUmfMPTP5LYs0U63q79m2
3sFFnO9x+zOp5n7/Ssk1k8FWqeZvz8LMXgbX7uz3pIgPeuoQ4sAnKIr2wI/xdn/6A8HX5V33kSdq
r518rodrlgew5TQGFRwY9iPlTPAMPLGFV+qj7XmmyFm0ifiBe753Q44zKzJ7vBAXtLStcsqUanhx
ZeGVwjT4EekOCHW6Je0tBxkqCIJHLPnQX+zgHQPho/Igf50voi+tCcitCjO8O+xBf8jHQBZWmwDo
0XohkW6JhuDJr9pJCi0pIMkDi0mpsCIrFszMSLq9AC6lvvOjzhJv3aEnWREGuOuHG+xGhzhlosJJ
OHQV174bPZtVPOWe47FAPE2a2fIPSIbHtuNqwFtyhlA5Jn1KIJrOpkZzcn+8ia/r9GKeVekHlS63
mkZ6unzDZOFZ3jYWlXxfT2TVLfcOSBXhACWa14FnOQCrC2Ej+aGHWHNrMOtsw7sKnrNZiH+eAW20
UnUyeitYEM2sFN3VqvSfgXqZMmtITUppvfL4CeWYuU5aUbApxCRTn6XCZg5kutbwKh9kvavSsDws
yDitAjDbDdHDL/LJhhyYp2l42sr1BNkmKT163h5xCDY9zOANGDaK8hJ8vh5BwiS4l39SYR0Y+OIT
v3wV1xynJ6Its1QP5EhmkM4i4fCIpyxHZgnR9MXLV9mCxa6koTm0g/99+bxfyDEGOJCCTF6Dm/Iu
JTL8UR2S61GYTWxvO3GophrUYRdNM5O0m4NqqGCKzXODrSCkv21hnH7rqJnvR6gAz1jvD7lLf7FA
ZlZYFEG3FaumkG4wbFppRrRiCUs3zgUEXwQGI6ughDiBahEVknwYF3oT65MUS3RfhlE7YJ409Su0
+zRnJF5IVRLtWjo7xgRml6V6rkW3XuUxhaCSydX0NVWiMPOmdI4IFEf7Zey0I+FhPKpYPeiqNHY8
NPydTmqvRx1FPUSnCyV24KQ97KgRJl9eMexkhiN3Dhie7x/SMP5gY/PsAAXE5ZDURsa34yKMrvR7
qcQe+byPV7eZLzvzj4H8ScW76nNXt66dKoZRn8qfvRRKPFXre2hpVeitYQmbGBlpNf5LQMxW4Bmq
2NI2EiCouqTD5A4/amx7hqhBA1GbtY9fB6WBkaYrImL+CFipYX5K/Vp9VH8sCTATc4Z0UZ/kETHU
6TsiP/Tne8LZSkb7lj9F7aNN+C+/q/ov48hsREh9K47mfOWhaHm6eS0knqlwkUFzPW4i0rcQRScz
eBuU1nNso09qRoxbiSVRjkkiEwL0APcL1+ygwBbNDOZbEFFlffktGOjf9AFOUxnu57fyU+mhYmNs
SnsxtiLggz4QuLC+emf4b9Dj5ue+CpdeHb5yoggjKhklhuULWyjDR+EC2CmRLtFLzoUdYV3gMV/W
4CIOD6Y7uDY/XBaq4GgEMTBnsgfYs6pMDgBsSzhO444mnEbffGE5FTZhQxFSQa75BBWr2MMDJfSI
Vvw2XAePFx2reFHghIq2glC9jTfdpGsLcoRaFwkpO2i1QxJvpJuoDsWNJWnxlR3OQF3g7kiq2+SS
L8T45JJaA1o2Fn3bYfKryZG7QJLUHy+nAQf52hwem6hRf+c0YSmhpVmc9fZcXJiSiDnxOm6jiH7N
/lGFfXa5vnMj17n9HPTRAIkoP4659ovm3wNk2eiPx8Tjulh/yOW1IJGjy0t1dNxxbmVr4eSygB37
VzObiuZrPlDZ/e1VYlNv7/16Folk6qRwnC/KEq+zhW0ydw/+JfCQxkOkWGtlFeo9EPsr/PVL2kZw
YdyIuYLTsBi0rrhQHfC5XNQxZ68Ed+Xh4QmOFid8dgY6447W9XJ/pIdoFHi9nRn7UcDjq60PacKp
X2fzJpFSdJGQ4Rdz5Ko9j8lX6h/4x+Akn7rUk8e5Saw2Rglb3JsvumoW+ZjnNgtp62GN/2avRCkf
4xlQ41DZVJ3QpVTqBA2H5X1lONbRgcQ2mWb2Qunrg+1OMBlgAwYw91i4qpBtSH40B55Qxy2F4DOh
5kYrbCzvTue6ozsXk9gC/B973uEU4H7zCNquwxqCskmqsnu/miGPEfTrV5CrlptUvfnlZitv5lVi
uIrWiq1guHEI+qox+zLoOoawid7hmN3RKIpBolcIwf1LDOYUHmtOcZh2egDaSsZ2/wKjpzk8dXne
VMPO/A4xdjbyMk0/JC6CJvsQUKRjqaahaiUtjwPJ8UX6yIzM5u3K+dWyxr4ODeQaTXc/W4e4PfhI
J0Y+1v0PuBtfLXvvg3e8XGitdXXLi3ZPd/PfgFV3WPo35F6AJampbVK3rGtUADceksRByY8AOjOA
xrRR0BExuZ3tgMS+9I+y3z2RPZ7Y/qMaTkYn/OPoINfXDIviN1gJ8NOE3ji8S/AmYuQP0BaEBPBE
9LWpfPQTZYuIrLwpKQeqZ90TNoujxkAgIMzjlm/ULFb+ZYTejn0IGPBiAanCcmydoQaNF2hTtNtw
Zuqa4Bx82Ld4r0qzRPOXSawpCsxSS3CrQYbtDyOKhrBsP7a45uRG0+na5spPk91kwQy4IpvTfMOv
7hLSH0oYG1+0KFWTo2JrO4p+KNe2MICVxsA3I4IqCgF5kGDhpGVpW6pxA8Yq7BrLuMhTpxOX/vvp
2sioF/kfc4/0ZzJKF922BAmeZ6ZZ1P5/NK9m7KWg70R2ywjjBrzcqf6rvhIiHH7pB0Z9SKpwgoZZ
rH9YmjEamiAfdWkHXR/Wv80qV4mnCTWuO5rgV8oMVpuUMTjAdX+DMGVoBel2y3Mxrqk/tB2l7aTV
OE5NshQ6ctXeZqstBwwbFMECXiVF+zvSoXxLLSVmTkUD6mngTCgzEYMSsex8oKhlzK4I6TUa/IHP
W8d5TKFeRwRfDZHuBwE5C7xfo4wTTplW0JOFrZQpUqStuFK2bfIMX5Zlm9++HsRPRvPtWKspFsOK
f9RCqxRDIPoyn3MQo+JBG9AjhBqPRvpZl91yhrwEVSWu/wcYz3+zvdME9fqaoqjcc4KJUQdloO3g
gso7LkG63daaz7ui7znOLevV8gnR1ciA7ckgg5Wd4N8ukekeiljG4mQkFzLjanzgn6o3pv2DisML
9qSwDLqjIptZTrohVGF7J/UVcbOsWurZ4Kf875w1liajc9JiZ34HDV2M50UKll/q6UzC9ATHZ5Ya
Z9+xGzj+hXH++FGJY4Ji7LUdsKc49xkucHvGIJ0utLAHjxn6hW9QltxjRlEuS7XunX4IU7CJx+Fp
9BD3Ol8cpVpMK7OfyLo3zJGWtCB+RtHOp+x9dlmrHvxJx4ljrVVaBqxdTA4Eig0JJ5wYT8VsCxUV
GyAv5TIXb4UucMOLLqCOfx3WOlV1XcJ5+oq/OTnjLlKEIU9y0aPbjVEx4NYVkcOBCu1lpnJ3Bup4
cHXZmxJg6uhP5jdBO4YGvHqbTo3OiqN5wykLc/lO5/3YcU/RRSA1BLHYbzHdX1V87cd1wkLSQufk
JdAZv3xHQIh2ZBg6UcOT4J245CSWB8r1rTMEUXbhbMT3TRxenTOnIc+URQNReVzWaq7vQObX+Sfh
1sf/ObMkh+1BTNU0t1xT7U9AnaD42aEqDcCxzH5LG6EmebQxRJghv7/7MHr+6NFcZKXqVsIj+IQb
V2IsqjrWGwG01bAQQygjlcGVujNa+zJQl2lzRuq+4LHOVkaE0FA81Fxda7a3APS8ALgF4uR3Ur7a
7Zh5gY/NfMaxlREiu4K3iZ0pVlci2HjR++q89AF9nX79d7FFDI07SQRqkKjjUSFkCiB4np5yty0+
F9nOc+cByWnTGFrNyri0w/AuzwApw4QKW4H1FeplqJ0XQojYIvIn1tdbu2A93IjIWyEKJz68y1Kj
svaVQ1Keh8KWul9iDxoo0Bw8Z4KCd2WHGPESW4CRI7P/4EaS9D0nj3WMrpLXhGkhQRFmo3MSRN6E
0s8bn0F8hyiE7pSVbSMEj6lzMSex2YsmEsnPrKOdAqTK7kOIcugviyBPwkK2ccOZ0baRmckGF9Ra
7FrREEVJc46v7gmvb0kPTVgjHKQYn7Jx22PY9HVxT8bhDZspgUIdKhuab0zr4Fr5uE5nmS8LIA7V
9LDE+xpE+Gpul5N4n+DpIfbskVsxKgUT22Q+fPx+qfS7n2HjMPbCb1KHGarT3WyfUl5jDEZw9Pn1
kPamnk0Bcq3W4rZbVexLUi7vKF0awo2DRbWAmu49nE1XCS/1dne7Sdxg+ly9BpQqyiL5A1ZaQtWo
w0bdYInLYHiX2J2p+iEdCb5M0iSrcJmxQPDmM7+03ortydbwSUp3PrsuTbobIdQA+jp7loHRoiuL
EzM4LrrkWnB4eeeSxTIMKVPLJ+xQZKfID5KEXxnJsVSRemoXU9GZ1wKCVxIWlOwWPDK9pL3EmYQQ
a7mHhMlzy4DDaTSij7RcDZIpUD745fk2+CN+0FP5vhv3yPKdfHb5vM/xurZEmhEklfYmVDMybw4F
5jvk15pWfXswAp0/0ioFVT6gwhbqzwNSxI4ZRQ+StJIPLclHrn/1PKcDwVADvtLNBhv8dXydJzqR
QFmOxiix/uFgmNAOklzwf2Bj4QABE2NrANMWKEySD6RxecKaXe7hpJ85k39m7b0wy3pvC7lEdbbj
yM5SCwUtvONDa/vLkrupvIGkQERetqTYYH9OZ9Kifuoeukzj7vAteU0tPmrAyIhHXg7rf9XuVGzj
4dfF3V4naGqVXF+Elo2y5kTyx4iybqcUgiC/yaaGPN6Hjrr9KGIB6jbQwZR5pjaGVRaZ1EqNz9ti
M9WVnalmiHtipRv0u057pKITHk5GzOW0hvOdZWz+YkASM8Nn15PJ0Qriqz3Ib2sRbouP5PQxFD6x
Sjwk0W80qViLBm/iOn40l8ftMH+ucsEFlPtyZ7+ybuNu61y2GFCg7c88AXZrBXOcCrQ5dUdXBjXd
514shevO8RGgQpQ6WzHUNgaJbvYuMSK5xCRUYlYofwvWdGU3hAhJzujQll3iLAHjF4BPzqt+N2Z3
fJduIk/UIUqMxCseA10QSzMmIYOZIcVYM7NmGTL3PQctY8nH3BtvufjJkvJwswEENmXeWd9FTGAz
qto3lcQwQq3ZzBbKOjdzAPr9JrPrJ85fKxSSv2Dk3OVBZ9Wb2iKVPmmev4BAFSz2lOU8rPyzauyY
b7iSQuSoP4KX56z8/dgVibyCDJvBi/2OZypmAu1Thx56kooTC8jf2DOxavRKoNcg79rGuvZsBuIB
tiTYsweTZqnoQVju1I0HH2uYLcilscfN4tQ8OrL37UF1Ug6yuYaW0px5r9+STynnu87h2pPXLLvE
kvH5hLyDNEXaAx9m5X8k+gwRuPNMKVHjNqe1+w2UJWU7kzOWiWd0q5dn5hIXSTujPJTH2sq4XQla
76oSrOolxici+ykT5XQdH1cWXlO5mhfdvkb2/6u5a/kdG0HPL676y/0iDq9N/ZI3CwZ3H8xiT4J8
sOm7fR96VsKyIt0mKhm5cousg0vvZ4XKS8oGbTtw6K+aAixc2Ipnm01WSgxhvjSFkj2tX06rpNHM
ViXhqaSPBZYe9MUE0vHv78kBC5WQ5aAm2ksvGpaZOmUXgAMzMzrh2V9UZe0qY2Y4UCMhp2QFM9ut
bTkjEx6fYhm8XrjTutRTzcioLBuqS+Ao157qBaeIdps1NzR78ggNkatXKEbwa3rAEwzGYkkbRfQd
jkhzQbbwuu/Hilo8em7O+yVu82KfzaVFD3b/SbcuKKCrzHCCgjcfZPPal9t2HZz5E3xXGfVaMnWF
RcfjM2kcMIWJ6s+shiA0ikJQLR/k2LmdUnREySmGmrIHQRZoNMIY9m+PXxwWdYX8D6VhpK9PIxxs
U7yJaLEPyyM7OYyqfp2qhLzEktZdztv/+Hqdn7qQZvOFmaO2gvJkWV9lm8oIjS1V7kzNoKW/lv5E
qiKl8PBiuGG27R1AOReFNadpXbDmf8NpL4jW2NGOT9CJS2IH4S3IHPIVfr2ECuGaJ6eUthxX9HmU
qVRtHNi+ZEx+BotjxUKvxztxqNifaOxemHoA3YcxqxXnDt1PyEeoOQ7dM+GLeAcJvU4tS8bjG72F
qBT0XvZFIGPq1+cmIxiRvxi9EVRXemrCE3gjOsvarN7z8LTZvHY3suJvsqqE7vEYB/Zi1cuVTr5d
22mtl38WNM8P1Qgn3eEcTVc/Rqnwws1ldejT5UVSzVYlwVMzvPAczO5EYCLm6OTPn4yuXsPXJzqy
tkmGL5OmEQTZRa9ZAipKmzoAYER7lF4lkUc+4Qca0Ip1IMUgfT/m91LYAfIxHp3GfE6s5WGymD1o
g+fIJfFmCUp5BO4D03NqDUEDPlnpWaXEI0+JxYRUc0dALZEQXaGqa9GbyLgVIt78t70nwUw12c8F
uB2XgKEEo7p9HWg+dKSOO/6SaVhRnYWC8NUrhcs3TAmqneI6ZLdQ3e01Afe0JUj7xytMPtGqY/U0
vAyN2F0HkmM8zuB+eFK5J1a460P1KZsIl6jAOJOELsSN4dWtqLcxsbkYbmC3m74dHalM7bvKNePo
FqoWAoW5nVvQc4yEOk1WGCY7kX3d8AgW/5smeDwcC+tsyW2AXohUB9k+i9MeMpnAmpK+EEZY8ihg
lsWcENn8JEro16dFGJwGgMPfXoqnp1Pma7sxUU6xZ0YVH9P1v50e0U4LRrZ78xR0HjU1zEIcKLZS
NgQgdE0ZG3UxaP6xIItqlCZ3zxyNzaNqB/P9k0P8RQSjyEBI14KIs09PrRdf0K5wjScJu00oMgBk
eo+/UB5AYsFzEAGXBNY4OW4+vyNc2NCjC1RRT/yNmQgVq26kTaW7oOHsl1r2EH+G/B7rSxTjSI1D
gYBYkhVGrSAHM5Uxgw6itz8Ak2e6tfi1y8/qXE+caJ38alUmOvQ8sIPVd3a0XWTHuRs2u5FH7Cge
xQyD55uIAoRaO3Hysozq8gz4iQRvLcPL61uJVvn3Ur6KeCBQB/eLX2OtHGzsnuMSSFTkuzK/WQI2
HYPmL4X82batZcCm3zTT0YFkTFDTBzbaKlM5o85TDtGK64WUIheLDRXNxgGQP1DKSgMQyLVKC1et
o6TxU+msetzNm79Lo5aep2uPIthdfdGPEG2ssHtH8N3E0ubvtMpylXsAxch9Ub/ESby4rea88rRW
LA5hRf7cm3ZCVTrKLN/e1gRB6Q4s2GANxjEeRL3eEgLcc/TSXU0gqmN3mixVpg/JZeqp260Hztlp
dNt3bauIUV0TaprPTJ17dGN4C4hVe0OBhS8oZ2ZD8YcVqqz8/D7FHMq/1B+ZNTlp2fymQMUmQ0Iv
JIjRgxqHaT4NytvzuDpWnGcHEKSWX4MV7rfetR2FXrfrvDu7CP3vQhFp5RaXD6l3yTgzvDquRjpJ
UrXuphuxPr5+kydpbAWOu27dNUvRmeRrWy7Mbze5d+rHX+VLMcy44OSVf/BTx8sVNmrYjP2t4ZX0
U7WakKxFW1SDsglTNsNddP5aZbfdZYg9MJ32NNnQHZNXbB5iPGWOHNbdVGNe1XySufZhTzzm1XY+
/pu2Q1Kald23uCT/4/QIztZ1cLTCF/nnB8GqYWgQHE4N8SpCw4v+opz4XnZpIIFIPEQgV/zAo1/Z
TsvzZzymTm2ss2PZrx2ZvIlncY/wB3ZD5wygXNKrK4ioPB98kPpBV/7U5zS0DWTw4vRnK9iBlpbl
nmkAgB+A+i2ypiDhhwVcHpWDJo6hnMxH3OjWGK2G6zAc+eJQOICh+3N6eRi4cvjICzZpoFJ/HV6v
T+GeArTrElJNCZJ14hFEVoO8wLp5QKNnxDYqku/0UYGzDJuCT3gD6r5elf52aw3DWKc3qYO+59K2
xSyQi4NmhuBKZD+Ar3EXMUa8YZ5OCGDf7kg8kXdTXJ3ZmJVtTUEehbx2Pg+8gcK60r0mo/P8iKFd
V76DeWt+kR2vzvgF+L/1aeJ6gqfWgE11fWVffj/oaN4pN/CACfJnCxT3E6GGVUTbeKGmaVAubUdE
Db7ARbr/zlrbIo94lycKrB5rDTy8z10/P30ugxkPosM7CVtEqMENlNt8apbwPFjMli+CIRrSkPNp
qlSZGIQ7bjRwSBCkWvSeBv5QlGUaPv4dVTH/e35LxW3TGH/ZlgatY/lYu3xUFO+zZApZQOeYctTu
6pZZkJ8A5GLeap+E165HZz/J2Fyk0W865G4AWTHg5ufWa338V53bOXkcRi1qnEuS23gbHzz/BFBs
jR9awsy9ZowS712J4RR+urfqfq2iJ9070KnYbhUJcgp4yEX5zuhyqxwM4Y4LU5IvbYTRu6631oIt
vAN2ZHJzhBlv2M9wq3NkpMl7y1thBERn/TMqC29PGLGZoGXwnXvuu9sjhLkgQCZhl2L+7iLu4D03
QQiVv0rrFEnrVsXUkD5OLMHwJRYuA9rzHc010HxiGrgfPiShU1GGk0OTI9mkbaYh4TSQleiKSJro
PyAN0Z5EFlYMv/OHQFaQwE+0FZmmUJ51h0WcFsd7ENhXcd659oFyIqJE3L3l0aMzD3SeLxEBArmn
/LKSjV5H0a9rNgbBu28aAarWxFSrGxCq0rj8rriXIKy5BKBsYzJ2xat2aWVJAtNsAVRSydtVeoub
Rz17J3tMZL+1w3G0ht0jlJ98QGPI2YzCqHUPj93vPviHi/0RDSnbML5+m4hAbytW0CWgyiklHvsD
Jifn+EoPzXm8zgFJgv2omKAVknHmb0gTvZc6JdubXLONqTAyB8kcDqU9SRLeWqXlH6sWDEDE808H
csCGmeYTGKGpoo/ujBZxZ+58akQTV50ZeZR9gbPLetc8u0NGQ6ciCXMtUwu2NFkh2a1mKFzREOVx
ICeTiRCSseAtlbt/pylSTJFOFeoOAcUwNAr09yyFGGOH7RswdxeBeqPJJWYHyaJA4A/UPjX6bi4Z
jkrGAe+PkyhqGIZ0jeIzFz/ldW9uKQ3Bnk4uyzjbArN05SaEw8GBtqnppaj+4i++JXOq3Z6V+1ds
3oMe2XiKO/nBX4IEXwsJGZUo1VnW+akGnrcCrKNKgNL84V8d+nrkWXsdMfjLuNCkznDKSdMRrvnC
dFEOS2WYv7DmIPd4+ISFJhz2tC+TtQuyCE123trgTsYE5qd7uUk4WHSbrOkVDQTeZO+qSWqUU2hn
aaX3Yti6OmrLvrinPLwoc3FIet/L6PfyW22PuKFrM1+XXqcneD+HTY2Ph/ow5AS4YX9pN7n2TX+9
cknsrQOZbgvhUxciQ/MhLpgZrq6pEK0ubuEuyDuG4U9HCd/TfId4nhBPr23d8JVp1fGNT0IfHjsH
WT1gHlvJsKSwvd73j3WnPsLQJexUzXLPkm5ooqBX8njT9QTVteJNbnpwMFv0vAcijacbK4Ksgqel
O3t/7oKfR88ifwINqH4NGwfU3ZLC/WtE50606I0hFjaP6wOvO2Ez3ccz+CJkKwYc9vRokeERsiky
mjhrn18s+EcK/eJEsQS3+eGiiPp5HY6A+bLRSYeZyVPixXhY6bW2cDPxnfsdvLeVA1ZPhhSbq/7T
TOAoc5+yuztEeihp+4Zi64NVF0OSoNIGuZNBAVcWx8ePelrOLmowBl8zq7xJn9qg9ohNdCdfyKJy
/bctDfDbioYaQZe0QdTNv/FS5nzTOZlicmeWL+5NxbVnYPD33lPP1jb4dBLYsPU/O/y0Snm8E9vg
JmLvgyy73QsNBEx4RIa9AeIdA4YLZvPibeFyUw7yiBGDl/od9gK2C7/tC/Ra1dQu5AQvzT8TC6VN
7FuHknmrv5UGAyrJnn2vrbYDsQpXVYcUT70XdQUbTVdsBY6imlLlCCTmslM1b0KKCb2Pp6zKea/y
J/swjkNzB/UNSwQaHpKKswcLtU2HLRe2Jm070Ign42LsPFbMbvaa+Pq+LxlhqOLIbjx2v0eXr+za
NtFmd3xJhXVUzKOMEX79rU0tbT0N4AtxVIuflpJZ4JY0Sa1MsCyFSgOPL2iC6Di6AN5n+LUMCqtd
dWBUKLABI2+y49LvtXRjpuciQCJGdiqwMWJkSJQfEdkHNpowaLuHSHqUC2BMoXAhYekzB/K0OTfB
wHvLXKekTh2ME1E8xK1ovL19lc6DoaoaRdOslfYilv3BLlsGVhwKT0xO+opstu49ZWRMlp51NnEp
SrhU5Le68HlqMgFkNbRvTs5HnU5+qBZV7bwbd3RQBGjM0QD118TVNWSe6YF43AQrQy7Jt35WPF1n
/JhM0nbLPjgZf4TjUh3mGaGFafmZVtboRST1JMMBWiMycy0MG29wLOQvJF7gbdLHFeXTRzf7Idkc
zdhTbGGJhyei4qG80wL3KbYPnvPX15cFPVf0EaU4kjZxzFX9AaPd51N9Cdwp9+mA7MgJ52OaTjNC
6+eCoUguQ4QOAvUsalntg/VQGb0cNixdvyUBkeFNoFR269QqurE0+qeOTupTzaccl2Xku6AJ0/lq
1/Fbp0p+qPGVqzSZ93Xi+OJNXpEl8LTPoUqp37oJNjcrgPFnJSuIxGR08e8vIZtNZ09OBXA9KlmH
IIq+zd8D6BuQaRIyY+QZdaYaPutPi6ZyiLks552y1A354Z7XZfXxpJ73XXAWPIHj2eiAyvh3QMon
tfUQOxZ/8xHzNdashQPaWQ69l5ZCT1L9FPyjtmtdlgoqho0u9ORrzTamu5Lp8JmFdgJneOMFNzfl
lNwcYDDu/Bjx8EhwM7eHZi3dwi5NkiUwbJWETvt8y1b/dcd1gCjsWbsdfiTfVEKSGP9+vBYmPiaF
zN50ygz9SdyQQIsS8oZfFG+YoJScrAjX0jMuJ3V+2gnS/olwSL/CReBmDdImq8S7vMU/XRE6zQtN
cxRBk+dm6c3rhCyNSpOq07+svNGtzAU635soWj7pqFPT1/TFCMJlt4wZoR5cp1KBp6c3aRmIDcTR
iMw4abLcatJPPTvcqOuLqed5aXFStKTH90Y/pl9/eZdAoc+wy0Firjv/ooM45VNL2c77AkKizTQr
Lz6iUj9LEeZx6qZEa8TGCgBooYTwI/BhjK2kjpPBnquSrpcvkMkgHDjX6Txwaprk8NbEVosimnSs
JGB/Q4B3OARMTJZNkRhUo9olq2M+CntulBP0SNool1LAgE96QaX3Ye/NKDEpdnpBcVD7PQdx1gGk
2PIb70Kwa+oE3ZRVXxm5ks/vtZbyusO/12edmWyWQEKi0ggCSHFWlhnRyqJ79oXmjHv7Nht/Pbj2
v3y8JWPNYBBsfHy9EFoL5EoCPTWSQm6W12uuuSrwTIuZuPJtcFlPoDY1wl1R6t+2SEUN8IUdVH44
3AI5cs0luZEqrpenTd5D2Mfzs6di/YoqwtEr+Ma1gkz64zBnoKSOuDgSX1+7l8VLmHbMfSZjJvaf
SY3dN0URX29ZwDfsdEwfahGuaZZufwjEUGQsRns9I49kcuEYj/61CntlNqU12IP1IWgf4+fHBLoq
7HH2/ZiFP+esaZfj3dIu/PHBqjQHKCv9hWcKuhRNclnLoIvMzc1lFwXAluUNWcKmzg1/M/q2ScqG
zVOeGghnW7C146pmC7TExZse8Ar4SJxL6iMgmDkUNr/CooJ/a73oGBdDuB1M/vL641+qIjwu72Fs
gj/mMFS/qEAuo9lSiJCUcnIjRNcJr0t4AeCcXR3rQxK61C9gXlpaIK23b2RyChUMn8A0ltn3NiEW
eM0mstNx20Sos4cwtS0fmujYmH+lZer2kk4pERQkdePWp2ePVcllmCdbkzcKo1JEStAHvPSaIuSL
IwSpq6nuYdhO2pzth249sk1fdfB/YoKRAY4ukKv2oE+pE1+wPXzaR+6eFlkC0LxYqaTTr5WE0+N6
UfQIr/Q2gwvhCAmDlV9UERY+VQkZlx9iOPxTMR9SNa8aESW4jif/GcdtJaSjuG7Kp067jmOt+e79
3C6uDOUfavx3Nl843hvljAINkk3i6vG8xmfQ2KrG4RorB1Yhpn4H6K/tYpczmHTVA4IWYyRXmG5B
eG5NkcPHG58+Q0cBnAzhNIF45mcCvuIA/3Surm74fh7jIu881ZjykSeJEqx5CGnOt1f0ppS0skL1
VcvA1Awj2lc7DdcHLVuvgOZfjy0Q+7/labHpunQ2EAZAGGCUJqA26oBYN6QO5cVfxHpc/exPy3GM
9IODRWGfPxYqx1PnZr8A9RjLfm4ArwkUnmsZPH+Uw7+OaVKy3AIqiZIQvw36xm7ME1gBBqCeqvq5
aRnBNtywbfYl5kaPqgg/vB/D7qB62ZrQtLEPpadLJV1CGSKE6cpy7+okf3XELtrrOrX7QSWaBRRT
1LXmFVok4AO+GwIHitoiuS1pd0WYcwFZmJ1s9HW7Ksb3VMb6uq3kjl85/6m/G4v+KmqeWj4IYeEQ
dB5VTT0rKNyonehmG8/sLG77cOMtrTD+je4uw8SRD/ooIMgRkwQd1HN6DA9fG8f+nugkb5RzOXkv
oyiY/TzV/ZMGChPoo6q3mIcevkouQecePFegyvWip0LDgT5MgA6MRd0JvpsWwOfFln0+FOvrZZPC
KKmfOppgwHhjsNeCswNs5tCFihVp5qdpK9BSQb89c/kBK03Yr0799DU17pjVOenLv90HCHf8W6mn
vUNJIW3yQh3GgMpwx5sADA1BCV4fXr5EL/g2oHIktpPbmb5Lzt7DCdgfRI++4rm19Y5zCovlYXdF
GMGKjZOHmnENcCLHSp7vUjDcKqLpHX5xapoon3lv3E7dPFlSrP4aVW/b27hQAssWUo/zr/zCodP6
2hpqYMslFh0W6685aWqSp2WUbenFuM9iCExveZzGftK6UPUziNLamVPNjWAlAPT8GB7ZTABq1gus
EHmdQdJOD1o4xyZFsqT/KHFW/92J0h8ruMzIRSa82eb5L7UOmega+ZsRw5rzioeABslcY4srAeST
WcN9EtEy9yArTf77luxotb9XTn5naIv6VYeREZveq8kBr4rHzD8DLY2/Z0Ejyptj6pfyURJyXjbh
4BuWZtk0zM66vj+BvRozglfy3zY/iVs1aiLcfFv1h4c9KmJr4Lx6mxTy/XeDATgrl49uTnQbcSaD
e2F8veDVU0PJ1bD3as9H+pZT71z+o9yLLyrRZXGaOL/oFcHF/URYo8BoF8m/WmeQsI28KGaAeIGT
Gzh8U/tahXOEEC0uyknhv/ez/M9peEUauwOZG8f8TTZsM7ChdcVNYT6vJSML9y5E7CV5V5nh2Mri
b1jg3h+G4Mx7otct7qAA13SY2vxH4frjiMj74WZl8nyvnUK7huAgMByYqeIfjE7NPC3r8YjEA0Vs
lQLMrhoK5nIjIeu90lrmpuUFOOgPA57ermNy2RbJNbOWsAYNYDqMO3ZRnendWQ+d7aXtZaxCTTdP
fzFfGaiiGiLn/BumSyCHxxsNI3zFRbvhkAfeswdVcmFefmPeVSsaBdAOgSQv86P6MHIo5Q5Pmcjl
G6M428jblokf4Dryqt9BlwOopaObFvxRuQurr2b5GLRR5KL3kJPo3/S9Fnax3nO+RyDKiMzxwKTL
MHlZ2R01zSNJtPKIZp7xhdWaODaK5nPwxBnCHExSrM6pBC+sJnOiVYAhKPUAoQQ5IWDpjekztcfU
qf/6gXsSnSJZNd34C3pAISCAG8OZ+o8uDhGORIK1nSKRM3b525Qxz2PRV6Ly1aFju6V+DBc5KBqQ
6q8PALF5x8Dz6bwE8y47dXMLRGjC5ecBc+BWfDs2RInMTlfrAkoaTjENPIOROe3ByvEV2gs3F+c4
VFzn9K0N5l3gpXOL82j/Hx9PelWB2AEM5EZbhBN8Zsh8CRk2jHRJ7rwnBe/AKayfHxBknO3u8XG3
9QNCcLOykryir+D387jnTq2pAms3qBhaeBXBe2OP9izsnOdkKXVuRa24npPz3OgDrMLXGsMvM3oy
98uX2MBAyQ1Brv20rwr+eLYq7Dx9pDe9057yBacX02UQHAJEvZ5cr2C9mdSw0s22xrJr8dIajmCZ
Wzk1tk3FJUEmITAR/U/4Nbigeh/bes1qEh8LeCVX0QUmT+pJFtcBH40ojX1+KypfNL2AKQMkIwQk
8kbhrI7XFNJMTAWgK9SDssjdzCfBhT8EGm0lD0ZqdZ1xbIhZXKoMIMKGpFejgyP72F+DQLAc9q/v
+NLjBWBKdq0ieZitVrOpKGON0L8CNpgms7B/6rsWJiftypsdfzN372eWaXXZo8vSNuacj4qo73Xk
KELu/DKvMuDVR9xoU1J5MrCssGfBo8MeDPdQMBTqKlQDQiIyZZqfRn7zSlD9xAN7kD3hQrA4D8xj
sF8Q4nYdlFyICgjyl1wji19g3E2bUd6Q5saJniwVmcCPZlcXU6+gEIwMNPC8S42kxcanfSYDqK8P
HJz+ZqmJ8ULYjhetJHO3N96rgRJxALjy96q14I8vxfCh/yMh7iSAeybiGLGBE+3IsE7QDaofZZ3G
um4RcdINhnUZwI90uBz/LA3RAwcqZTx2zexzFX2LbPYS8M3Kc+z2MurPWhfbYCTlB1ZarlYFeLWO
SwxgeZ5JW+i59ZmIh57o1ml1ZgHXQeEUtiSrZUkEUDbgQerec/L2/43DLMZSX7+0tDclrmvR2YCw
wB135KSkKj06jLhaTJqhAMYDFHu3ngPoQyqDiPqdJlLahkrgadQZqK1ujGk8p3KAR2glIrZQeXxD
9jEqVuHjRni5ISuyKSuxLrc9/01s/K3kT4uRGc+xo3je1QQhY2gXYLrvR3PAnIIjFUxwh9s6/O/Y
K5OCdphgDZk4eOUsyjsl8yWyqik6wRPAkyyK2bKxIghD8m4q60aOhfJaJp3dYhtyrakEYLV2pVIL
s8cuxeZJI2hZdvGGCiNfE+/XWJheWN7s2mr/UpuSS4StT3Gcsj4+6xd8aeMKJquB+bwWJFoGE5JO
RNumycZKsmYY7zMEH/ZFY6rhB6U8BHsGGlt8n2Esast/dK3X0LArFeZ57ERkScxfhhGztqH+Z95f
a0V+FjahMwzxH0nepUIOC+zd7Fatf/zMSj8IqJOcuJFPmOWUWJK2+Ij335T8ehEdKChaXDo/rV1p
aVJXghr89W41pEDPhzDWsBYDrH0HMPwjhfVr/x2uj4zeMHIz92P1pnPqtDBl/Nkwzxz5mPkXjYwN
SoUeDdB6HfRLZ5N55jciHU/xnuYwRWATPAtd0Ge/Q4wDvAJe3O/O4b8wevRfmfLvHlQ00SHMDZNd
l/kxkpY9nQ5KPPoZ+k82E9lYao/fj6DJ2jzv9XzQk8dL7nDODYIQ1GX9APaY6/WVfauuJ7pLojU2
SiG6PiTCnz6qEDU2a+u26VppO16gkxgxUtXxFRwqupzoGdDDHpzXwv9Lw1YdiIdlcaeXJV7a3nyl
K8/SEO03YjbbFW2zidFmfYnGjmvWs238Qspgqh0VaM8iYTc3Y00HxfnmRYwkFJxzpt7KlEtLa4F/
roMkmXF+mOFDbbL8sD0SO9Rw9VMN11j/Br79TAS1uQul8mH8ze8Tg0eeu8mV95Tqg92/kMXg83Xy
OPqw6Q2OCesr05q3aOka02l/SMLOwKsD5qRiJFleFgo1lEEttKz3uoEYVWhRWDNL3FF/tXiDE40q
mWlce3Km1RDvQLDPuwAae3WM1/N51jRvhneAOf0PczZqftohYAvqB5jo38RBIBb2WpvRYUHtfTCl
ohMxKU1FQV/9zgfRPM2FtaggPhqoNGRC/Ra2p3OgqdzLSMfpjXCNi3vgsQHUmJRMSFy+g5GQyjOR
gDRT+ZBD0b3qfUo8iOBToGdope9PeczBD9AlCc4O4HJrUPv0v+4ZcYSx9lYzwUMFVzUydIuz8+m6
92deovj2Ph1jxVyTx6GpDX6o2x4Uj+EKyySr2V583U+tIcHq/EMCKHQFWL1//thkm4dg/SVpN51V
quGNOjgu4pdVXEOguAEUaUuqamU7f76RZ4zWZKVyiivVry/uYqHtJW8RKoSRq/kDbiUWueKGMuQ0
O08F9rogOigCcIUkYZeM0jqf5kvgCcmjC8tybzyYvM+/QCS3dyIjARZwxrFWtbdvCGzw8k0E6cxW
x9fduk1osdHblzfzZejShCxaYYvvkkZoEa9lsJQsELCW4w1oBBC9SL0NWwT0psyvzUyiHKkUtPTL
EocdPKkMNg8xIGhTSMn/fU55Wdo4RyKyk3J2ZHDeEXeSvzOCEeDnALa6i/vz0gJEmI4MF/9cLQD2
ibrEbpbtUAw9RAVlp7gNRRiBp080gLodwPL65xJbYi9RenVmA8aPtQvRK5GBOGMB4Saw9Qr9sBN5
fQA5ujuofjqG97Y8erE4bMnUU6x+r1E+IEULnYGQ5L9f0LZ0oKGQuc9y611wWdcs3NQtktesuBFh
IoKvNDZ/fowZ8xifgZZ7Gq1iMmKeEaNdZkx5d2S8n9O64arYt+4tYnuNiMGb8VTMq3MBy70sNY56
sHpKuj47bligMRwf/8AdIU8CVFS7sQL70HnsdJxkQ1vsno8J9sMM/HJw/LSggLBUw+uC60xCPeJa
m4EvEf+jkg1nrlNVJ67GIf0fUScdNQH90+7ixqnlzRG6mQWr4jVoED7GmA0YdSzpboqLXizVneiG
SW7/PZNyivl4Be8ywD4Q0iST4MfTf2DmDAAEmBBiiK+kqwDb1cpscSyt4mEVhBZEDWQ3iFSKCWb6
cGMhMVNV/GGv/PzAv/cFMe94jx7Wb4T6m6mspbAsQ3DOBBp7zGBRU9PPd630BVC34wWuk/UxGvQH
5MAALSKf0ywaFKbcxy1GCb8KpXGI6tvtHQHt9APM0G3bibxTbYKTcz06AgmZs4Rsru6PQO2hmpL/
0H4zAxqw7VVNRoIroB8VXvhX71da0Ucy5wwExhJFD8aCqiqklwfv4tWkOTy4AxONtL4xkAJfgaRE
vvlLKr/TQBTIqVhrhIeUXMjKjvk9q8k4D/HpIxK3Loglg3D5Qom5TXCJHXWOa3FxyP77azfIs8uv
hHGw+AU0RAOJAyfm2mYmUvpYAoq23uJ9hxCGCjC++O7eFz2FdFf3e+8sQqdA4QoIIDJz4XNnZbpw
sV2qk5KOqONV03FfgBvX38vhMpuckeDc8L0NC7r0MS53CSQ9n1DMEdrKr1D6nOTS0lVWAh2D9bmt
eXkUa5mHQR9y1sAnQNked/y+IpvI7S0MPQ32rncNR3/SNLC34jz3LFSoDFaOZ2Bs+iHdF8HNHSr1
f4XfxIQu5dmYvQ+MUgLEW5OZzmjHYqfVgGiclKmLp+CBqPV+zMhyGLyVvullKMkX2Q7KAXuE+s+e
2cz3WKXbxI/3yNuD1Vabv6HMrC5qWgCRjaqqch6ZyUrQkYBe0kOiUDYhFbR/3q47Td6VRugc9mzJ
yzjPsXdK3iBpRFOLZOMVaM8MW4Q0J/EJukjg/NieIE5F3zkgCMIBuOXFSdSjb8v+HkkIgIsqds2P
f1Gs9CYrXP+vkoRUxcQx961i0I4CrwLgbbFWz86Gvg7a8cgWxRoE/J9WWIo/GoadiUTdBiWEsVtg
xnFHJQEoR9pVi4a+VX3XkxJetBdO+5oH7gEqz+3CZ0zO4IZfNRs8ec7JeA/MJJ9BjUmw5cfAMu+7
ox/T8RoyS48CkbiGdhs0DVAR3tj7BhTurzLa3QIsoUPELpILWVC54I2C39SOkCueHgMs/7fbZHsH
k00Mn1z+9nGFGgvMyw20Nr2wHZZV7YhDz9mYjynIrTHfvEAMGuXitdN4Y3SlOMcwuVovp89kCxgy
M7/bsjy6u6I1Z1D64w174BKM59Hpowwtbb2kiwFs9Pm3AVj63GMVjlvOfOFcE4BWpOizyFYP8IW8
mSEYqeNnnmuDM4knO9pzUAQ/EfimRla0g7zASttvk2PExkkF5nVJTx5FUbTqwD69L3rRDJtUXaKO
k1ABqICdZV6Uc6SQzxttQ0A3XLpL9sb5qg6wpH56+pGN7gTiNkfTp5bOOfVWZKv54FhFqKNjhWLu
0klqEvibVQFxXJb9W58Y7gCK8L6MV/wiurIWWq20sX0sdug+qTRKD5cytDEUFp11xQ9gzkBqYH92
EZy2k4y6lRwEo4yrBnBVtematef3QTkueG8L32/L32yiaXpxA2w4ei1xkCXaczEyM+Pk7mQSM7H1
f3ALUXYtsX+/nsqBkQwHFShza3r7dmTzOe2WCKIfjC9HaMqlILYgmfVTLqRu9bvNk6nFdsa8LuQ8
kAZJr2JD0s/rDnpyJCd8pu7qoI2gMgOwfsgyVFh5rUG4GbAldcRaM9o4h+iDJRTv/th+t4dI82rS
YEb9/W6KPGLZo8GKa3juz0BAHGsOBOa7vL0/xQe8uUAs/pw9fdR8hQZtiJR06SCC5oTR2VzIu+q8
nq6lxUH/YbLWYIscXVACEEs8HbnncgHVYnG6FUBryykuXf7y1R0eBuXgE+nrqwfON3TF/qQGbCIc
ehJXNe8R4Ag2REXS6TD22UvS5c1ZRVppIf6d76h+Sm2vZrC7bShW4orGvslOafOAmU+wDUMc2KVY
MRe2NGQGQK9oogQlCGGpmoCa4lM4Ya7+EDzsJUnb2h1czGw7ZcjS0d09npOWYxE1rbpteIJVj32b
ecOoCY2Vn2IJfUOhT00SxROKqfRtYCL9sBYSgMpjvl3Hxd0b3Y9y33btqJDiubc8awhmg25UaLgz
aP3DJQdf0MmCBvAPIZrwlb0Oy6sntAfweKgka0EjhgVYvaMdb5GEgl36p8z2rmBhuqWP07juuiiz
EMgYFwTUeABvktfbq2ddy+p+X72YCUPZIAKRgltjQgeShSLkoqBy2ys708hm0n7pa+CmLBsAXWzT
L8HPvCUuoN7M9tl8tjaqYbAhyT/esS9vxKuEz8znpxIi+6VWLnL2kTh6j7APj9ypeePIcPqP7/kI
gZpo+WM++d0oEQgGiyIeqBNeq+pA2SyMYYdOya34dIQgwTzjljszXgGKeFl1x7zQCnmSlyP/76Sz
Z/h5c3h3ZG6s+CTcoeNRAdtoXhw5BjkTx4bzKlSbqDBS3GtNJ9hxl7Hi2Sf7tsKkB62wGcNivBlB
mUwKGqLyxqJUMe1Hp8xzI5mvrcjeO56kzgHtgU32MhhOB/bJnqxLOkODJ6mufW6Jrz+2StvnQhDd
IY8JN1uREJ/j37EIIkH03gjMuav6qMJcVUH+4Fd4TJ6bBWgZy6iCdAsDEV4ronio6+qxtaCUCy7l
NGhAm6yNkMD9SvQaoCSQ1GZUOlUXbskAkA0iQjyRC+zt/kkFg3ex2QvU9OiUqCLVhqOxzOcP4H3+
dvJVbeVu2fXdrQvQXwwmFYKZyAmDjEJPKnosFzhLz4iBgLsFZioRDw/Segv19pTxICOrY+eFzjDZ
a7l4YiKEE7pklvYofXAWlYys+TBky7F2xbRChG2S2XnWbIwEDhYAuJEGlZJzQX5YZasOfU00mOuJ
xRJD/0E5/Uvm1z8XDAitZ+SsL52yS2Ck0oFDv/4Qssm4fV4pcjuuMThyxsDOLvaF+00j946SLAYf
gI0Zk0gAvA3eC39vQ+pnPFccMnpKxaCI6jXHfR7pebgUjvefKffFb4DatBPGAbox0cc7PD5Pj8ad
ARBtJCS3JAR99t+Co7PAqrKzeB1FmYxgMwlj0Ha7Bp3HQkno5WhlYM9hDA0inMKspV1YHcgl1sYY
ojV5oO4fN5Swt7BMmoJXGNGLEjj8mYkQSDqU337YGH0JZ3GQds+fzHjxxowOO+2x6nDGPSmQfOSM
czkosVyQE8sMt1S2RvJN8W/BNgEkrYJh4W6/48qukqq4+8oqbRq2iK7usSJc1y8EhU5InJK8XOQk
ZOgPFtb1X1TglPLz/DH9nC+PMpTB8HMDYi0LCXJR4qJVRk8ocjy91LJGfeFhathru+v3MaFVFxgm
N4GCzvf8Ht644iz4uWEUSkpkDRTNcsvblGafk8p3B7ENG1N/kO2GC+FS3hZHGMF08vmk5WyuK41W
i7DCH93dCcQS4Gsl78Vhc6ejCldqJZa36ORBv+4SzOYVKIt9gR6DfqDEwQqNE/XlStG3cGMRUEjr
AqLxyZPXSMXxhh5rKb33QPajd2URFyY8mAQVJX1p6utVOw0ySLBJGxriCSF6GczjvgiGxV8s7Sby
7h/+wX/WtfkGtSawaA9eFJn7V1ibwGt1DedWNAYeyRnWjIFguhFPIM6XZW1J1+RKR0FSK6mxJiJ1
WYy6+gh5IOpXQ3kBINMnsQIEsoFL/JfJGqFuDooCCR8SRb+LEIqdAzkrqd0P1jH2QIRANR831Kn2
uIv4Fqw72QSELy8vlV6NwEfZQ1rTWggzMCTKrmirDosmO1JnYeCEZk9iHudk2Pov1gY+tdyohztN
poFukgKBkIgLpTuyxYjq3XO/hACL3Gl8UQoUlPNl4pOoQuNqJvQSySjDVY2xkUv6cggPkrxUjozL
qWK9bK4+kSocr0G4W5lUTwYRl5eS5sPHylz1ohHye5M5vY6yLPM1b+ft6WEolMxX/y+8X5yexYDA
joXa1zI5XyBOpGwdwepQRRtJj5R+HkVmLrm5DDcYIqTMJ1hrT33brz/cE9Ka19uC3DPR4vE/gBiv
1Ui/0UOkJPe/Utoa4M3/jrP9km3Db4It4Ara7d+0zh2XdRzUDzNSXhPI0y3jZfGnPYFq2L8AB5uY
JoYRiosMefflDgwcZG1QDzPArFG/0sfJ73sUzGCpcYdkhBlGGFpqm3t9pJb4oGEnAFTB9z3cEnv3
Z+82IOwFREcivuc7J1fhrSG+tZlmmXPfg6f/DctkzFfuzGKursiV5FQ73qOehXzE3TJrJILuWvet
04SOTXFUx5N/n7JBf74z9AsXNW26sD2ykMNcF7fqcTlq13V4+cpZV2aziEwoDqZtBOJ/DbWBiYno
EjJA3LADxdgQCW0EzZb+QAY8FOm9CAv2L/ynEJT/zbrGSnnmesGcMO+ENdaeQ9I7IotTH6Jbt2Y1
6FYsuNOIoCBFHi52UOFuiaZOlc8GIbFNvQHwY2LkqBiJVjtpbTgacyKcD3w/Tw0xmsPzLAQ5bL6n
ZXMQdSut3LkNtzTthYfhRMXPQRxKhs7VlH3qMqGDW49TT9G/tdnoTUkotzLN5aZEfgmrp1uyceYz
xRO6rZRGgQH7i0KykJ2UzrXlQ9ABsqLtd74EZn9NF81O7Z8Fq0ML53AqTYvAjXSSXs0CNwaMB7bD
/mq/zwjODLrEqrXxlfRX9BbLJhxPnNZhZoB3dQ9wPIUQK/tLYOF98niMpcgCqJGHAxNU6a70fU64
Ep3oWsnpHupSFcTJGiybhDDBCSEt68C0FiqWv2wqBf4r0uDzMb+/+55pmkoQJ2rZhyMiyxeDzYPY
0g1VY15+b/xh7oU25KMFpfXU+CrlXifPcPJoJBpel4JgEieiC9qiEn6VGFFQabCL1NnehQQNMCFB
j/fD3Z1DrmuMwK2pOSOPJx8tuPaltZRYJ3MgTO94GpA6UfQ5hiXXmbZXeMEYhuPDhSZ4Aa3Croz7
HGc8XEJYAcJlZaLS2LgNm5ZL3UdBkcB1ASHUShndmJRIRcQfo6NICrByjddE4Imc1CyfCZQlXyRE
wfQtgEQg/zYMHmE9BFbjvr0tbFb5n21C8aqlnR/P4IhN8cBaO8shFODuKcRmEkctNytYzQRezClE
4i8Amck0qwWaWZl5klENZmXGohTYew8nP3LQDy3qYtrr/QKX8sbd8D0nve0nMRtaANFjzfMPuuwU
DIlu4a5ZGLQ6zWVWoQJjPaIMOQ4mz2Dm6N4Ebh7N34HlDfwF47806zZB8hLn71xFvLuSDGfuh2tV
aCykB42L4d07a9l4fqPxc+hCkMfkAnLW4Pj5dryjQtdICwEsmUUaj8Kx/t+pZiD0OWby3MIwO3v9
r+Iq+oPGb7B8Dum9P4rADwzC/UwjWH8fU8/iKkJR5o2uj6aDizt9WlmT6blIG0QXBNVEJaMqQlJb
dCV6G2N8L+tVs2KScXgdiT1sSCF2CHp8Sjwd1e9rj2xxGWEPfFQreqnwLgVAH5w1KbL5MrQmVq7m
eerh4d1C02hpjNz0cBs5rIlI8tF4vOefxojtpvOmdWjrF5Q3vznrLzokL9A7eyTwOVF1kFCCIcNk
E9JF/oq/MNiKaeK4vsgEv0w2aIpH4JhEOPCsGZuNeq9NSb+EcTIBXyhWRWIsBLENEPQDhvYsEqma
KQAnNK91e7rwk09SbJFOKOxOzYTNL/t/QcSoW2i1VXDgKOrHxIWOZVUbc9rty5ymDgE4EycQ0oPk
Xna6+NhuMK7yZBpB0ML6P72mDAvijnkbmb+UFvIfqPOMExbFE0K8dDXLflWOGp4yEWIntC3XiOL/
tueIiBWe8B+hsSDZ1xjd7Ur2c0RtCUH6Vc01kCVhAlNbKouRzqEsrqjPx45rlnwc5KbfWswKrzIk
wLPCdKLw6AeGYL0AK2odHyeFawg6BhyEuTnthl0L3iV1i7SUGNUGROG/iLDRFM8adwHgsuWJFocp
UDSpQmQ6hzK9dLfNw8JpQvGxCaMfreo94MkshYlKPiG/zO1OHYEHBikUwNHYTfABVlisfEpekJH8
Ll5v9sM6LTYmenzVV6+1Ptpz9/ifdFEeYHn1ahm1eMMjZQ2da4N7Rw1m2cAHnaJeVn4mjV8OLmkd
5LHxh+im5jJGhnG6N2QgY1MF09y8BkF9ipShrfrKEUl2WcwtdM/pIpsoLwIaFM/fNdj6CLllDsUM
vtwCLuOYpniLacs6ouOEp6zhwyV2ihgHRlwcCAkegnm8RMDjoIJY5DsoAOk9f+6vFotUEwlxfna4
pNHKP2QX+98i1dDVNIjcJeXGo7y63HEZdTeVvDUh2mD+lyacb5H3B1OeBxFBiBOUCUw1metVM4LU
eI1a+mEa68qP/6ElxGdTiKPfMLlzJc8E6OIMs1IOYSiQKgIFcL/6bm+m9T75YpzKCghLb8weRbR/
Z9WXUsL5f4TtaAgNfQvwRZVeNyfr1/30Hg1ds/UEsOfedE7uzYqGb0OjZKzHiN63+FaBQlfHqg2s
988KVAkYg6fA5RbR5uBupnZBuSPgjxjUh1nVdIdERMhVs7iZBHHZvG7pRi/cP0OXMIJmniuh0O3Z
fe6IZ48ZNe0p3IG3xD8/rQsata7gf2o9DIXpSnXuw7DjEYxh2aATtWhH4SXPlZsittKrijg8lKd5
Djh54e+5AxlBO0d1T6NDollEX/33quLvYCfGuDS6IlUnDXMUBg6Dn94ldCC+ksQyzqr3txrnBZs5
OmDmp+7Fp72xGVSoalcAgO6iWgr2bfwKvAMQc9o48nN0j3zL9VFUH9/MagT9OlN3vDB0IqmcfnBz
R4he5Iaj8AqjUwBgWONPcmUID8YCCq9NsZ/RUZJM+sVjoi1nofboZ21OmLnU9uYbAPcyrd8zXcG9
mZfsvxWqa75rYPD2qz9cNaMKVlz2vj88wEvjbM1Io9flbfxOJYduI94iKQhbI24+W14gdC3oikwo
HBCFVyF9UBBHw4U6xu+cVxq5V4jm4jU3mKnH2CQ0W2eK2Um5+2DC8oY3igDJFDAhJ8gCtPun3ONw
8CUKjVW3a3F3ZC4uk8EheJSKNAAnu7IHbQurhPZH4o/LAcBSC0oV1gUqz540ZT1WrIXZyt7iILfV
INkS/NCCQZC9qb+m2J/k1OP40nAl3VY+YdVcBtlXK13dYQP2UQfCEIxRIqRE4G5h5iNLP2T5HRsA
zsSKxilQHIQVCV7EnuZCg23tjV8kS1SFCpO8pWE2KyyXifDicligMel/6jEmgkjqCQ6TQVIPxcR9
qcglKnYZkj8lg/5sFOmhyM7n3qPt+yyZjlXfLTwrwj4QhZNGSBwdkIlXF0bvPnb22W+RYGIAbYAg
PbMKkCOyHGBRUwwnOTmC8usELQUXoXVYXI7b+tHXJYACPLUEMMIBTyXBJYICEZzmE/7P+XRR8ExA
43Ito9tDu7V56qGlT/evF/pTI/XDHpL2eBiVl6a3qYfkocWZ3efcoBA00zpTWNJn3uBbeCt2x8Qe
8Yw5bO1Xm60CvCxUZ2s4UeieyrOA0EhI43qUSLbPUNt5n92M5azgfBtvKUp46uiE/dAk9cBQFx6U
JtyBZHVy0SbqrM5DMMnoPHTRHdHmniViAVUGIA0NiSiegYO4gw7iK/JRMy114wVo4C0bD6U+JxDg
o9EOJMRaQxZw/dH9Lxfw+5OuImzy7qTw4CQ8F6rDm4VosuAsh5Iyf8wzCYdUFPcUePMGX68bmpuQ
U5JH5RFdEQ6P+hMWadpxoC27De/A3tsJm4zx89UxsgVqGfcx4Ravde9wkQulcqCrHcHo9QgmPYXk
fe6dKTkKH4h+tXoSdja0rHmaWhWIGrC7SEbQH5ik3xjrf+JpthJCZ6QEWjNvwNaJK6mLIAIsd2Bb
GyEX08Yl0jk8+gMAh7/IbBgF45ARJllHAr3lwjgPBupLsdZq+5WftCvsCcvxs0O1ZARHHocsUCEP
dq8nw7Zu/Qx0wHmuVE+0M/PjtDCbA+4qmQU9MJQMcGCwDeqa+s/pWSItb/P+/WMXczlQtUMe3g/9
Q9aKld+GhbrGpPTNqN8Rt9RhjOLv/9jjp13E2r7fTjIgF6FuPWbBh/E7QwaEAsbUCwsXgjDHk+EI
jNwm7Gie7BmHmB9c4WUEVkpGGKNt17FDfzaDf2GHDIsVv4iNDNbio8vHGAVOsetXijqReJq16psr
XwsIV2q9TpRZg72J6cJHg+T1lPjE6WyhckreOlD/OqwR17KysaJFreNv4M3vLQWdcBtQnh8csNlC
+Ks4zXv2o1kp7wyx3gQpmrWji65fCPUzBAI/PMufdV8alVlQyLw+XnBxvUaBHFxVKZkn8D1OzLJb
5n+Q7Ts2J+W6tGej5Z0AOE39O53Qq+2JQWKmLROedeDz4a7L+MkY/lPMOuDhNEXJGgcHywilu78d
xTO9IKPvW8vJhFluSsZL7HZd2deG/ewHruaSnobAG61jnKrOBRLOWJ4M50hOmvGeYszCTfV8eyEb
Zpc0Wck0m+uxG4az6lNf74yfYKNTqZgn6X11JUouSYQQExYNoZzYOx5QLecoxH7LLHr7RWh6joxE
kmG9qGMcKkvZ30Dlteqt72TAtUYDX2mPS0IhTRCSzAe54l4byzNa8MUSGfA089d4XFBrtOVDmVyw
ZjovywYkXTLD8z7yLN+6L5EI7kb49kWPh8OalYix6WuB/uvs4pOJ+n9oDTKOLQsvrX1LIzx8aPSP
motzXKA5ELLgW9mytJRV4XUD7WcBbk7syuz2vTIwZJqbqVVZln5bY2rO+Lg3zYJhw7IY/jZOznWY
XXj2GNj2oMpI30JzuxGAOaDzSteHv0cnn+idzSiAbMNJ9SkFk31rUJs67N8tleYvNUdL9fhwsUfP
oOeuT4xAsz06NPetehjkb+wsiYPorBE4MK+VImqwMbXHakHwB+lETxwsYZDnuU4lbo7zHv7PuoCp
UB5319Ak7XlhSwdLOgiboYgg6fF5eURg6Bt6EZ0GgGFpx+gOjTyxQquS8ami08Rc3EdIKES3azcx
NWmo73w7VctttGzixJqg0poBkKD7hh8dkerpo97wQgGhS5cxErcAkMWZJm6y2NEbNQbGDwLtUBuf
rJ+qpQGA2P9ZXfRy6MhRzjnXzo4CaNaiA79bUplaS199hMYrlPFAQnlZt4AMSvzrvzSfgBr0hcMl
08hxMbiKj1xeOmI+irnepVcDd1jDOoQWmoEn+2COCS7H2X1wHiBVP3QFCyySl6i4EzeToUuGhyHh
lqNaFcZTs06GaHcos15/bTsmg/nUZzbC/OgzemXNjdCJ+P4Yy0jzK2uqNWgsH36Bv1srMYE5VmgV
aA3IBqgboJ8TcjGvN1rCKwzoR7wol2OpYIUsldvgWiInnlSHPUkbBCNxVXKZqafezZHzpSDAkoZy
age4NzFM6xJzzgadQueDDdzJmwRTQDtSwnWkSBwZ1hSh073dZ5ykWOM/c/LAaQO9Fn2ZpQ1s7QnU
IrW03G0gSjP/PkEYZdioey4MfR5mltpmsc0TcR1jWByN/C7mSJIM5TSRTMiM6Z7Q3W2U7xyIEO5v
3oO4yVmqEJINfdIDUpF4CKNrsirUvCF/6cCOtccOwkJw/H1SadZL0vphAEeWSH8R7L/X+Od4BcIC
1kHSmaT5m9Ggd/yGLZq8UR9533V33xvl4sbuQtMSINCH+VxBzh+3aJ/QOBjcotx5wP91lev9EMDB
ivccEQczzkksIn+TUMBeY/VJ1sdPSY0B8CHwi3IjQbkQQzkNt8qyxk5F3FQn5KxScbsrmgdCMx01
fQjFPJuPAxFRNND9fCCwqQy+ZkIRcOwnvAlGT36TJrQiw2+pBqFDuzXYCGgaSfbX1Can4P4GwX+i
JlHYmYL0UDryUq2Np1lks1bcREXHAsHlVjYuncKgYMdQVo5Q9HVD6GXSZvxDJDSUiTDosYGFeKKn
tzmrFxBXl0+yoIrdbJERkBGnXcQOo8a/kQxzEH48OKZEtn8g5t49PpIfDg8UHg1WHNX6Ep0pq/Mj
EQ9TVXewEu5bE2BmU9NiQVA4fcVVbo6waA+XPsjuGO2SerDB6+LQExa/QKpIbAaGjQR2X0EqSN/N
ywbhvvB0evHB6VEj28RKYOBQwVBYNNz6XZdgUbA4Zde4Gia+2mribUxI2Pd+opyDuzb6TXyA/eNo
fxcvpjxrF8pFVxpMoXmbrwRnXFsvkOOmXwbT8fUvcjVbEAFfs6x0YiXMXz6/2mG2RhMGjZ66md4/
+goF9h9849wcN7vajwHsN24t9W+9lbhYhab4DJR/5QjHZLzON+VIUgomZBREQ19CT8IroNPNrI/S
X88eomeSDqpIS5KfC03oN5uYgcbfcj4uQ5kUN8XVZInJpTqLdQVWHetWHSNcyMPrmy9eVkGUSGr4
wOBaQ41eF3rbjK3LhfQXp13uNrIh/sdq3cny1ENBAYF5RHBgqBslGsbLXOjys5CJgKg3UgzJis9q
2+1XB3cTZyF7sFa0oXSeoH/SILAAyRsTiwplY8quU2wbjf/o2kgy9Fesgt6+FsHIZe1+z8uTUSnC
lZaPnX4fdJMUDwVQv/lIav/VFI1zHJsVVgcik0Vs9g9muhutHHktlgIipw4qym+nFhCI3BUeGi5L
rjOf4Fisn7EHmNaWVuPHOlDUu+owaaHUQCXTXywKHcHLVIWdxuhsKdtaiGI/k4ts6CNjnbyk9pay
RtVOgFbH5ZGp4xOkqbL5blHPGx8C7IhKPa2dYZlP2qFQ7Y/0hBPquhH64zKIyOG3NglBmqStxC9k
OWgj5zNGoead3dnOgTbMtCDp36DD9plzw4zn/aNq9wNk4Xn8/+W1EWjXKlgSOvd6NOEQ6Yz4t5jy
J27umrgr/FBQd2FynKlL537O5LWsKagVMwKyM7aROtIOa1HreUqUlYSoCJYq8VklLZwa1IwO7jDb
P2BgKplti1+DYT5+8sjq7kP8Ahf+uSuj6ugAmv+dp0XrDyCaaUsFd5l7HSUUPLCnjjlFdaPLTAWV
eud6RhIaBTi7x5nxOaFyfr6lR6QLigUHOs3DuCcKapfdlmwBRgwtEMxs8wvLe6D/y5WFBxQ2xnnK
crzQQfjHvYJxUekvSEKyMLKaav4ZMJwBduLTIxmDzPElSrFLaNtCBZGnUBccLiN31HO1QqtMjtDv
F/c+se8Z49IESIZhHywwT7PAaj3HZ0tdhRqxfjKK2hsn1YD5dY/qaP6IA7TKMxsZmVXzuHOGodgO
a7+grYPdLVR0eX4G9PpmE1E5zkFKbeVnlk4Db4IWE0oaPr3VH699k2lD3JTae8Pj7D6rBdirXLYZ
szPDl5JadIrL7k3FjwQjhtxNOEgalrdgyjlLB0R6vi2ucEUGZpnZwhLHWqgrQxLXuN6q2C6OrJAZ
crsLDTExqALe+UmpFk3j9xc6c0nXOA0N+h2qaPPo54l9dyMjhreMTtUvwj/f2DA8Mxr8H0MNqBdM
PhUUeoZbAkA6Ip2e9Df7hHEnB/VQ/x4aPkrln3jYHOFCZPlCCOEQmojQY/ABTAPtGCBiWWMGBtP8
2CHTez7e/yqo2QiUarpNewVlSdGTjILq1iOQKVp+WVoawOFNmOT+wR2sk5MnPLg6NnPolF7NnaVu
T2nHICeGTEOvqy0+pptnQBkfOLnmZpij5BQ8jYPtTJQHkYLvzQmFMuPGovLn5YHqsr5i8a5OYEXQ
2pyLdDHDP75VLhSh0/hy0ylOtNjLlD41izl0/zB5fIW4InUoQKblaejF6TRyMuj5TmnvgxelMiOd
HO2FNNQamdjmBcoQfWiAKk8OQSwW85liKlN1Sr+W6Qe6bE+4B4xq1lBNR0MI/zSdF8jLCGMV2RS+
RXT1e+Ivea9xv9s/214YpN8qnBj2MpMLMlGlSd7KD/wDy9TXCLUNm83ty9cdiaG/FLVOo8o3i8fC
lg2Y/I2Qf9bz1xq9bIcweRbvrt1ufxUWVNWMf3BalnIWqKWzdt9w8KHHSfvrmk039k9h1pPabsSq
cn/CC/2Bp6StJ09/JMueMa2LWnDJQ+0qTA0+zU3DU8KYWcD/NrNL
`protect end_protected
