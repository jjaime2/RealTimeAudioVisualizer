-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tUKk83ggatyrJaSvicJzT3xm/gJ61+wdDhfcaKXVM8ayaWYGcXLVYnUYcAdg/5LER4fhyVqx7QsE
KJm1wrrJU6EX6tQEqVeGAdGVaGbdU9K4TJIk+evppfYrq3bP2ahHBVrkXFSOj1OkzXKUGuMxHNon
Ou7MUAxEytK5BMWpLUEwK3dDDsd4BaskxEdYvH9Cm20ta0IIheA/RyagkjpfWsCYewSw0BEU2PjA
CwKi0C1LRxe41cjPpTz2qXhYks2i12GiXcRzPQIUisrTPUzbTvo6NaTevW5ADc2yDk2RWGx3zt+R
VUVMgymRS0i9/VhPBtJ56sOEj9n+8/uLmKeA9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5168)
`protect data_block
QT0e9oMdP7AyeqZKD0mxtBiiAnJcCJ5uftAq3r/SWUmmQazC4bxg4JNd7KzUP39ncQ59azG7Msyv
MPeeZthYTcrKHVufZZV79SANH86YkwpzBVmIG8FNSeOOC8I73CUV+XSpFlHhM3wIezFAbHjoV4a1
PZit3aUcILkaozB51Y5oCnUWvmF6KpfAtQaAaFeHMj9eaTfhoomq/jMjMAu7XdyKe0sSc5wY+EOM
IIGpj+E13R1wArTndjNMY3yMXs7UnwV/otLvTA9WnHa0e3S3OM2RPtxozbWf75JKyCnVJ4wP7hK7
XzZuAAfp/jJU/9ksi7UeBvK427PvRUGiR3gMSHyNGX2hp2EY2URGpHdyX652KrZRSmNLhXCM3iF7
lqoBdNo2p5FZ+e5VWKhoIUy6rdyIoA+pv6D2QGljSQPuboLIR3giJm+k0hABf7QV342GM1B3sIZb
P40Fum/ES7YtgwZr7zuP/Z/mjr92QE8WRb4LiNJXKjBYDG7MeeU4eMGj0eDvOT6Uj+SiLAD+QdqT
ItukGH03l84oc+aV7ZTjPcfwMy6XeGTLU1HBBk2DwojM4vuxPvY7j+7mQ8194hUl/Jxuso/+TBuZ
xSbs/AyNLlm/ert9yrLBYxwwAt6t8FOBgHDgkPzyNBxbeagNjaDABkVOaI2j2pcsyYpO5rOtRc2p
NiyrbugQLe5K9wO39L58BY7DH4GscsmPocGKUapnCw3dDVlVrSu7V+gt0pKt3LcYKxxvbtMrJ4Pp
+1IObVeO3Jk0tgVoAE+j766cnP06zRvac9EPz0wAiLhDpdrxpRcnH6Gyt1ATy/+I9lM+PNmUjzHK
/Zst94RVaP6jw4mYChZ3N1/q9LApTeaaON6q+PNYhYk9btD8YCXIK5r8QYEAk+VvuF0v/v7+Mo3a
Y40WmCcIh0zDx/aKE0b6b4+4IwLYBZuMZVnpVu024+DrXfZe0yv05vQwGQ6E74ciOWOlZGb07thC
EhkgbgMCWX+3oWE+SZ/91GL4MXIVA7IHmVd4aq4RfIGx0Gj3ePfkNYy8ZHmDhqSY/1CVJo5zF031
i/7NBT/1x3RvnuaXHanifycNq1jfZPwtHvGjIRRIBWWZ2l1EwyLsBK5Pvnc3ytJ6JoVE4hyvB7W4
L7RMITR7n/x3GixNoO2wL6tmk2tWiRARk3j8MbyyKYR7Ivt88C9QP+kyq6/SdFONtTEciiK3Prek
gi0c/5fm77Yl1fPUZLcLEGD1Vz6pd7248O9mATmFO/w/3Qm7TY5WPpeLk9CQIN+0/meQwJhDlvO2
UGChHNGm0cNeZ/O+43QG2dYLdEgRajKRjBTRM7d5zJetcc/MT2IgEYXEOr8Z7IlRz4f1MEPsAqkJ
jyR/4Kua/VfQX7L0WKwQzRpHKW8VOEU0yy6jkzu11JB7SPKqCLhdrUz0OBGVzmhmsR1kuUbg3Kvd
KVM/eSDub++35CfBWj3sWkffeAhDCe5qRbzL9V2CUTYYzK5qn5WNVK73icBRMnrTzGiE5lAO3blh
WvyTQLuARLVW+7ZPdAkSB5X1PLAvsarOATZziKm4DwnV4AxfG8ihn6a2PwoJEEW8bTgV+6ou9xSz
xPPHX6JyQw4kVzQo3n6H1gZUaILFb/pCjH55O5ZI4eKQh8g/hh7VUyZ9cKpXRhnDmC45D7OVHwZc
y6/AZ6BnhesK4Kl2pIoKJ0IS0X3FM+q7Okr4M0HlshX4LTtQj78TUz3zxM0dJbBki9Jy2FZ/6U8b
WBD6H5Wmw8jwKdi7mbGxHCH0gtTSF275ogjw0mWUQjFPHnHHKUWpDka6NZ6iSHolxAYLp4ZTcc9C
BiuTMnL+IjdWLVBraZc1v5f9iWWFZP5U1C4FlzkC+AjWWrjXKMoYRnpM8fevkNZcXmbPWyrxo+14
ynBddTfNGHogzG3+cRlw7hfBBvLvlVQ6K0A+ALg+0ZJTtlE66/KX+mXla6cNSP26RrUY3wkhs9ZW
VpE2rFIsG+Q+DcfBXvS6WTCfPeBa59i3AXxyWtHhmY3lJ2G72sAmtSkQQ8jVE9EucX/Xw1zuOwV3
9rmz2Ud2SUDCK1QPSPB58+YKUAPPTQoWhVEuqk1hFXcryX2NRbXqauRXkBHy4/P8Lw3i9oq8bTMg
IDUjX3JSmXm7OjIWQL+bNOr4X7zE3KOLQ98Zd5lCNM/GvasSNPjh2jf5JI5cHC3dF2SG76d+15eN
a3SpFWm+npgYQv9ymQJUnLawDSTcVnvVCV+HZfJz9nunX5EXS63G8p2fJsjo9CKnjyQGFZKsYfjf
8iSgoR8NFNAYqt4Zs3D5Q1uZJjK4YOAG8fjoyKUnH6FwFIvv3g1cTRFHtiPtCDSs/CZLmtsAzcye
ezdWpzwkPWXigcW5nTGoKfr5i9oE+BvbHK3EjXHJ9H9YEPjUhIvEbuN2hgnLQ8rEtuztLHOOuFUU
JRX9QYNwpj04zvlc1OUJNqoGZEwjUug+We7Zh+anbVj6j2fan5Y7wExU/zJ9e53/cTuJ/l/Dapq2
GtzIZMu93zGoqOmDBbVwIoyt/d8t30k0PxhQmR/X4RAAIRAoqdmK0TncbqHKdNJ2NEERRHwbffwk
SWWqqmnD5GqigF4vmzBbGbfNzwvZZyA2GYcbfpe0k32CaRV8BRqImMhAkFNa5YNwWK0dP+KbdTb6
Uvxfn+zmXmPCJelpKtV50eyUUwJqjVz6mwWHTk6lx+zLjq/ep+5XIgtV9rN1iec2VCytdsfHZBjO
ZdoVzz9tPTlx/RIZZ12IesulNQZnLkNEcEjC3kG7G9FY4ZN9Zpzov4/2gPPPibk8VQijJzHWc5xY
K+YYOP87H5cWI+gHXXzmZOzIqIS2qp8XuW/yEDHv8rg9F9JB2ZVoL3oNmK7gIOMWOP+tOxDa14jm
ltq6DLpwZex0PbokewaRu59cgGU//iwA4ld/uUXFaZNRVL011lPxVhA4HPRY0q2q3lFqzBVR6yHF
PvHC2JG36E38nyDeZWJFnzRuZKOdh1oIZxxT4DoSJBovVy0ZB/d95O57l/+bq0po/ujgMH4fMezT
gfFrt5pmOnPdmKShQOAHPOiGkVlZ1xgApE3UYSpTdn1+p4xb9BPzubKFR6DHvCGZbZp4vuojDOo+
JrSmtceI3p4uBivJNxRwrp4Pd7OJnJYic4kJwHV3PCuiWiqvNVYUKHFvAquzqPDs29y/8a/cnfkW
IGaFtEwvJWdTqvAD6jthoB45GI6BpcJ/fl5vimY2WYBwoPPOSBcDkdnn+DNHmHu8RWcCp5JUaVJS
TFo2XYI2WlHDAswnlmqF+p6SrNC4hA5/nH+0zuFy2zeepSOlKVZ+dhVJ4dErd5ZFVuPKeJ2KbaA0
hDNQ2aYO3sPHbs5NuEmrIt6vvM3UvyYy45ywWEs4G5bpJYbxHBwL4QR7YjCFbzqU0r4ERE1KOhSt
+RmoVmfwQNnAOz6GnSRYvZDTS4nKf9OGfGe+r7lNZCVt1tLJJ57rbb5gyVv4TZlbh5kk3lBhZIbn
6CTTGBJGHJY9+KErXfBKn0FPX0WXe52f1iVCoWLq2UpHYZrA8APlBAENvX6D2ljwxs+DvNg/xvkR
HaW6WyQ4c7HinqgAb9SXKKzZ/D7FNVLqm7EREJEjzSxMpY+R0rHF3pZDkc+LstEgazB3UfS+t03U
EIw2UluNoCJxtuNAr/ar5vg/2SSMNdcvIbe19NWfJW1wHVR5l+mw/TVDi8rCnAidq9Gs16I61BqT
ND6RwphG2xWFOSjLIQO6BN7gVpLAVkg7knMDEPIjngCMpOFC9cTq8edFNDkhDyNeXWZBI0i2/ksz
y3uUYA8pd+EK8sJTQ2bUCqwKwoBehUX16bmSVwKvMBAcF+WSQ2wpZ4U4qNou01WrzRFF0SvAJarC
xl3CH4PXKNB/M1zlBs/NZIPf/cyhxgsomPV1LpWhU3ndtoO0HtDBmPlp6qgjXoneVqArxM2TOZ1m
X3NRh2lSjFEfVRfuGaWJ/shc9LuUqYUwn5YPLBujNwv5LoNDmg3jJSBLtVwHxrtT9F7SBPBx8ShF
g9hVE+HlwRyn/DBgBRR9vg7yfLzteyVJnwzKH8psXL+/JoG65rrpbAeYFudMbRadu0uCKf8+1g32
FqLcVqD/e0EjTNwoQL+VGsUDKI0/NkAyCAMJ2/uTnH29YnyGSjjo3r/LUFbDMlLpy1C03+vlTX+O
7rM358GsAkAFxc9Fyku5ujilk+NH+5uXpm1eHzOuESe7TvS0CyddLIqhRF0+n2FcF5sDH9HVwU8h
0o9tWx9ByS7WLZCd7R72IRCjG0DtF3itPodmv4LeAKCssZmrGlnClwx9vdOBs9gBtwToGyK3/APc
yFKx5KD6wqGCd1SvjUwAmXfhAuAOYRGnO5Dr4ZoLStO58xRRp2P9bNFlN7uwKIUonW1X8AtNK6Cc
tvc/3PJXCMH9EG+eQEvUzeDVf2a/4nzyRY5HTP2J1BpGoCnMBACpqJStM0XsHRJhiaV+QeGQG6vG
at2b7DNNxZRMlSLIO9xWFwCDHrNa2UdnzmrDeO6HTuYKj4epY81UYj4d7fQqJkkXPqjMoCrTO8/L
RgfUqYpv74t7ITJ7I3+1UfCUSBVrLlyN75KQAl47IgklQSLreQ7rRIhKCj883WxXSje49aqRS47S
x6tzIsTJR2GCTW9R5EznMM3t0sI+V0LHZ/gvuyeyfhCsUMclWTBvAulmoWjASNPYwooBP8oa8rcf
vya5ZY7M8ZVHxSU5IHVqyns7lutW3N/4mQ139prZ8Ze3E5F4YiePugWqm5npzlVCDeTbLTBpYClq
cRDpD1qi1PACIpGdebBryEYJ+IDpanr0kYCaJ8HaRgaFz3CGdTcFyqCpDz0evMDthsgRQ1/lzbfX
ifseTWoNCPs2mwzrL0isfi1RH1gqjHMj8m8/aHYAswhLX9y3dPiqApr07+bCNOgO/GRR39MwnHZX
uHJKyeggShjbc+x9pasN2xqNlXSQsfFP39LWgr7J3CRKcFiKjyCvqLBMpXpewWv7D3cLiLpavYso
n9vOZRT93QpJx25gtEwAgAGWK03zMMl3V9VHr7hlXZCVGsDBmeVRRqZ3dgp3dw56gVvDsYDWStuI
xJzp2uHviYl4kWux6VUfecpFTKjSdj3TfnjQZSYW+h8BdMkVDv33h6SyWFVssBw0KypXHCromYsH
iJI/C9OvyVTJsOGRn1EyYt7dG//xLsJyaKihssdbUg4xDpQGBVBnlSczbe6i4pHrmx8xtJcUVlus
/S00Tx7+FvSL8K6dMwSa4xBVQeZ1XX0l3Wv6CoqilInFMhEx2j/xX36Hiq+wNhlVTQdpGgPNVSaM
kPspTlCtYEC+2udfcKCjIQrH6wtm0ss94RtLWlr/Ko387r2WZwU0vC4HPTyPprJes5RVR1ru8GBv
zOBCg8r3Hjos25qhQONBfIdpugn0JF61u63mCVIgfYJVtsxbFx4X5EpFi/Yey9XjhAjFqnmC8fzi
ow8rwDviSPXFk/kfCKMNUuZjllVaFNaOxNVy70E4Dw8v8TTkwg6yJc5IlIDpvAu36ZVMiIBf0toE
/hKJErX9ianTmypaUJxUf+R54U8AUyeKjL54VEVpzjLvDr5XqZkPqqQBmV1SldNyLNJ/8ngTUMWV
kVtK/Udw7F0lBS8CqY7Fbb41PNn/8Cp8ZE16JoQuzmoMYdu6Vq/BXvXu9A5bp4A5+69EPlMWhAyq
mR8o9S6o/fEfi0EndpB7qTCXPxJ9+93hHwl1ClPc80TOmZxXPKyxpCtEx77ipifxodS9LGwHU3pe
NIz66k+Pc1k2TqeG3ZLR/6Hw0iBO62w9ca5MGg98XsD3c9VYYOsIR9Rtp3dj/iXHMskEq4dWVKSO
Ftj5F2u4POLMfP+cl2NkF6iUJ7SHNugb9Erybnu5JOA+3KHUB/eTuGWRRpK1ziA2kR/p5FNKJMWk
xrIhGzJykZXSlKHSDv9s35KTrQl2J21mGjDnhtz71XW4DQgV1hCSIkqdo8FGoJ7LuzrBlWzOGQHG
0/wc2iji/Sa2kppqCNwYTYhB8R0iZu93sMYT2+jdmnpWRJCXTLmvcGoj5iDUwWShY+8tCk4ln4kx
AN0+EBRZfN4lpNcvBtn4D7v6jRTmfYFgOzhW2oo/o8AEt0hZpLJ3wBzCCI58GsjNe2RNVaT2crRo
cUKW2QFfTSeRumXmXsjWicEN9bADHzl8nGfO4SkDC1hkQiq3YrDzHriMOcf6sGpnr0r/XftyPxyZ
OdVZgWHMeVIDlx1VrUNUKontm4nD/zDVEYVck19Hk5N6w8w5oQ+E6zdaIgSbvO4iIX+DQDEa0MD9
9MkAwXLCYblKwQo9Z7aUK/C1OdpU0v8VaykD26wtK2c1SxX5v/VdekZCj88mx4cMNuxfLeJbjOAu
JXW0XlwXLhUnZcXdxLM0DcSO2jQZR7CxkcQGEWLfncJfjPOlM6xqop6QzBSG50fS5bF8rAULxmgu
rde9rXboFGehgevSnNANxT9FVnjpr1+d+gIB9okqUjbGYebQt7Ebqpbu/wYPDcUf9kAW1lZyNYeQ
ErBHsXuQD9XIH/sne9JZtvlrsCGwD3w1kP4VjyUdOWAC++D6uhCKKyfScVUDl414Sy2+Sb1pYB40
OQLz0O6huCPpfCEJgu2UZpnYAvp2dPn7tVLwGlqUO4/ReaH0pDp73JY8nZkh7ai5t5KRDwNolLr7
Njfn7nlqtytQgakA6JkLvuvxGj2WiMvgmHqhbYkmAijSywijKFh678lS1a1Rb74jkvhITkU1+ak+
RiyHUKLbeFObaNo14AFmjH7EEnPtOkIlPVdkeruE5wvZjlEU9VW4skrEF0BkyDg+hajhBYPJ12sO
1IuI5lYUa4lFT2V+1IIfSQ6MCxjpz7UfUTRG+Fdmd5Y9CxdEL4M=
`protect end_protected
