-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
B9pZScJGJLuaLZUGhBRJH1a5KgjmTbtCXbYsjz13EZlE6mExX099oCnxgnRn/SmQ/eLcFq3HpXum
74D4Q+v+hBTllFdOuvNvZWR7U5EOInvgVLnXPoOXJ74K/k+ZmntESdGfSFQ9q5HvHbd8eDO2czKZ
aWq5S+sl8DPWTLT5EvDi1Y8PFO9jmLOVx/aErqP69F0i2c/6U2SAoParuA8ee07VW9a/PjH0ofuE
PTk0eT5I3eytuDM1JBUn+rX1cA7mZ9h7nXBqJYcqNSXXqBjToBmzh1vtwfbnrXeFmjGVAO50qyNu
u6O0r22xf/ntOlX3dQ0mbJ+Ad9W47ktpqVG+7A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 83312)
`protect data_block
mO7YAAyuMpIiXSUQy8ExaNJcNC2fbxfl6k2fHmYDbleSZZvaEtqARopSU4G7XN3CGAYkLshHioxm
NrAhZi/HESACYtjBG1UKWU0mmh8wBNyvJZ0kadanhqY5BkcM8pWqaUqIZFlskRNQf04dG9ofWBZE
gil8f22fsXATEx2u2x0YlzZGAlGiL0LARlK7xOm3Zwkl2+4HjrqM4SvMb36aLqr6CfaYOE0wotni
fDEaiXEiHr3x2R1jPL3EfiBWJEIDnOX8IROcVZpyrUsAfNPWdbk+bD83uI9c93XhsMuv5VBL6bZ0
2B2r4XOUFsqD+PZjtG7KG4C0JchNP73iiid5vBgEENbxnj3QC1pBKIpTYjeFgsBOI/g2fqhlUp8v
oUjg//oq4FsuYU6oqqnJAyr554VTQhsF1/5ihlPjblAG/JZLSH/XwkAyifydI/Dd0AYE2lIHGfq8
oYfzNRR1yhyaJfyyT8hVhsE2wpEsvl7Dluvb+RVVIUDsYiflCiRNZSrMyeNExdIf5uH6IE4jazEA
1sRie4wa1H0DzAt29D0VKev1yIvNdnY8YprUnKKHMAu9cWpwgQr6nigS4X4IHBnil5rmoY68RUbH
jVSuIrmTO3NRnwx/pkuAqe/1e82o5M6rcNnx6ypFsXbI6WRosDB6dtwFnq/OwyCTo1Z6msKRWGCA
fZjo0/honkgFnSG2eADCsrpUOep9HfCJ8aanywStEReRziCA7pLATaRKohqG8yj3YOPGAacJ++1x
lzyjduV9Bc9XtTGJosmyE0fviPnGI9JcNm1ah4NlhDh5ar0SXbdNknZl6luMyI/hZ268xlelIvhc
/VZybpxNq1PKH80L3nLtPvUy2OB5aKjdFBNJvsP6eNmQkpFyckGqTmrjGgUBEeHThyXv1TsLooeA
XYIRN8W+b+EnVyDGiaEGtYBa/MgS12xRKOdyXmVvy7HdSuR9B4FLqvxhluVZanBTUqKlIEruaoMe
Km9Q6n+6728gDv8Ag4lkVVC7bLRnRqeIQAPbjo7Xq7v1++vK55y0a5iH/hbKUqyIySI+PxTTx37x
wnbO95+/Diozbn5x3jQvncHs/M8okd0oVwB1sE6eOhh8fiq988eOu1W+7QwvMfiZWer1o4EzE2YO
9zh7h0cJJyOTakyLjFtqMsOTMjAfrKbliw6JxjsB3I5upFV2mOAm4E3uyncuLM3CqXshnBjppuoM
u6kPaSgPXnpWI/P9RdSpDa1kjixKUHXpVfJxQmdFAzjzat751tJFngubNZ6sfZlbawiDz/97n4Mc
cn+9tp1+nA7snHRgMbIGIXDtRVhtfQXyqlae2rl2QvmbfbKn2SaP9rh/6XbBOH5q98Of4p+qIauJ
xWAiKzR2q4UtZy2IVud5PAtzLh3sRTLgzhTRQBcnBS34cP6j1MM6LCQm7WAP3hVh0Jpuo4UXTSxs
Ehuf+Es3BY0TXuHgh54hAVCqIz9RHYRnfSoT/1BGXJNld9Vus84Dj3Ll7CjzG0lAuRIeirBgKBaX
A6uRT9LaExeC0gleQKBZZ1nFAgWy431JRUzfK6PrS1nGoZ4jHYM3zWsb8Ux9SHooKi9+a4RgCOTX
nOM+NdK8Zao/FXkaLsOvZtjCBS+RkmNE4l8llj0uXWtKA9P4pd6EmnLtnhTC7K2AOIdQKNwGf6YS
ViqLlBHWw2vc0hgPeHZINq0p052qmGEgbffa6sDAowDTEdEaBT1Rq28X3K1/HNu4/LxrASGwlpje
bagd/myQ9F5gMfoM3GrYiiLAtVPNnjqRhDBP9qMEhK6yuGUbR4/3W8K4CfZrETufJ6wwk1dhV63z
BdYGnpX0cYihXPRKbHBX6XHL8oT4NN3qFfqu0IFf+czhO7oPgFfjMXWdaYkxlh/UuphyYp9jAyTC
AXbJZgUK/aMXZq21KhiNbgUMKSAdhCZw0sEUwbLO76cVVY9w8XlmnVDAglP07nq38+wdPlqbBNfL
lMR2zrxpet6rxmkjtpaCnEF1Zl8jw/76Kr7Z3HM6HI6zaDQuqcaDlJO4TXdtTXlXUF9tJuKkspOJ
y3D57UdRUmbj3jqaiGkefShWErhj1D0ie/QbQi9Xp3MgkoO0mldHT81UuWgbZwm3Hj3XQDrcwiH9
nv13f7MswIJLMJCqKDWAd/vIvKLx1STVip/Z+O5aYSbsaf1ypPc5F+D6NIWGZgQ4KLAuKs9k9bvN
EbhKKzEai0MuJ8YmzunOE/3o+Kdv7RTawEU2mVtgVlo95R6Yc9Aczf9ujrH6kVrv0bkm8mJ3G7KW
84wkxiTvxiyrJwsyVBFxOb+lNcQLCgkOddPq6fS/O+SQKmpUTVFyXWvN66swFhy3T77utGPSXrjF
TM9GQhOeYh7RQiz8Eexaw+EIi11P3BavK0GoTI+BwqR570RBihSRZGtLw+hMClEWpItPj340LuNy
/JdwITgco4rwmvgMurSO9tfLbEYSaJFEwruI5nAOEdZVEerzjFzGdDcKxiIh284JN65rQ0C4mP29
xxHYZ8oCGpsJ22jgRG+XqfsE5whprFjIGFw+jxFhI41tJGZ6MqfLuQQafiu4JyvYH8rKe8GshWGY
Qe2HlX1UpNfqeN/acfkrOYxv79HxlqUC6tzFP185Y9E4pd102hUEs3/IkUmCLcWrrjIAj72hRM2z
iG0VuV13z7DkmTWSoaEQzIOlq5S8qLiK1uoqkPJTXL29E58B62+n4OqNVg9KBn2OKgzeO7anRG4z
I/8OObyXzRYg8rmfgZlyLxMAE6JGqLqo3BI2dca+pBgbFt6OKdLQYdKZlXbr+f5IeKIee9HaymyC
FtyDQq4NAu8Ws2FqUZaHHDEZdzIhZq81MtQ0q0uE3elaYF4OB5tD6tYSaw6DiJIIe/SJFMCW5gzK
OuDSlyjCTaKIpJdAAcN1uYoLfdjapl5qXFuqOqpKn6gHL/EbUwGMjMzBr4t9hZma5tyFyD5xVJ66
7nipweNAcNtOTQ37pqQCT96BhrTOQopgmBTfa9XZjJJ0pxQCiDJXgEfh3YEvifpN9mmrbbQcON0G
XoWO46MFAtTQrcONkm9Df3XwHhagPdruwO1iKuuCBQP1yKdaK3ecBGRdTbi+chUB+u4HhbXeRs0U
EutqVgzPJw7MftFj77OVu8Ib6gaUfoUDjtiMBZ3wdoEr4zGKdtIyuSmEUsWBOAJWvXDFwa4q9+dV
g16i29wfoMcd+scHwXI3+ed1RcI/khB6utDLzXT1N/hv83erFiErQ/82aq9eREioCpxlDl3QK6t7
cHIG6J8+Mp+vSLyzQTdbkjl0diL3c+sVq5tiKVTLZhyLhyOnWTjb/aHp3zsfCPbRVPpiQMmNCXuU
wbfHH/y7wBKvpDqvjzi+1f9NmvfAPF7u9uJelb0T7gq75Oe6gak/ViFOI55WLIQELPmdJHoCa6M+
deFR7qWTCSAL/xVrqUlq/0KibMtOdnWh0/EEBX4Pw/lzG1w2qgUJHfBnobzhtDkGVXoaanBO4LeC
uqkPhDSmEgeFN/0w3TK3Zt5ACv1D7Pms2Lr2Rvh/zcbsRNK9K40ExWn++iIFmczTHVxutA9OedP3
ENeE1qhuR5+2o3Mn+t6CNL0SHEVGNtIuXMzWzP1Y9q8m5Gh8SQChbdi4KVaypPWdzhcSQ41sbvC/
jEAuz2idNxXFwJX2p2WRu83igkdC0M/p7dK/L4Ry2SW+Vk75HiqQYOvItdfgd/bKNMeUC/ne4DXL
6vEjwsgxtVW9QjOCEYFb8BXQpgXP7JGZsTfkaJXvrsxNuGnFOIIfh085iz2vMC/cxeya6NxKCPDF
1jkkr66X1z5KKH2009Wn7z2L93oL7rAbIfC6UvmMYrITUonBZpVINtiAiJ0txHiDJA10WB/ucV+l
yvhkFytRR23tb5zeNww3RLMy+qxoM3VRs3bfh91jT+UcSpXIUK41mnI3Fctga1AdN6lnjJ9jADeq
BPiOsoiuKLR1NIiwoXJ4cr+TKGRYfpp9dn0QUm5Pb4rTrQFIt3+SaLc9czFYLju/p0qeBqlygnVg
UiJPmcggQLK9DlIU6mKHaDqtk3VHIgDR8o5Tw1GwIFvo1TKP79R9j6uaW/0MWCTebCgRJIJ1SbUz
bTL0644GvUzv5t1NAPoVRjAucKxZ3SZ6VyKJWcdBSX4CgPGFUE16WNH26v5mgaMGCGew+zU3WYjd
jGFV023kcXTNpZzm+wV0VebBqEw3/s1nDQOxDudLqVozyrKYIXOAWmZUCXXU/lZRqkLOiuf7UZLI
+N6M58h5JIqFjIJ6SqwM2a8R6iu0aLbKOddioWYDJVOIgYmwI2s0VNALAFFtXOodj0apE3z+30eQ
M8O6bCYLEa5fJsZDwneaTfOsG/fAuZehe9ywP36i+/y8Aul9LKrA14FzR2oBHUXks6tj2jS4Sf8T
ZDejFg+fkUuXJUG7kgznxqYuKoTLuua43j1+7dEjNnwI1OyItYQSI5I7IESXFJO/AZwIxj0dIQ2F
XZ73yhFsRgqntv4vkhOEAyb9oo1uQf/n2M1NZZENClZHbhCu+8jq93JQiVRC1S5wQF8jLPnANxWw
I2W8krRPzQ247Lhtia/OWk0NtrvhAFAEAv0FC8qdqp/PsYSktbGfq3zrNYpeskMBsa1sQxcuNQHG
ku1wv1PU6gv/p8DeOVsl1sNAjD+ySdsxc9FX0bJIDRfO8P6t/R6ioUgt5EUGHGzM5n6OlWmvdK8O
rpyB6+DFkG+tr3Swiu0whGXSe4Zb8YdIkZCL303q9kD1tp9SDZHkhSXONzhI8EQFyDvb8Cu6gcgB
FkUwK/2sFGZGSb07FA7F5/ZINEp1ek9yAX6vLJWWfiJF/FPDmd7kLkDeATMO5xOC3EeC4yfYgxc/
Ijm/Rkgkpo9zVj3oVmzPhER4cApUc8qX3UioZWMixoM4rwXfZLXXG7KecQ5bVHtMv5mQ1Efgsw/V
RwmLcIZDWmgFy3IYwFEZNPXVJ7p4HI81YCcufLiqI0HCXgTpr/PfXJWNwgS+KbD3Z8CcGmPEth9c
/OPPovxYPJ2yjdziFAesnu4eXXcnEdpxUJvSwB7oLAMREsWrDDz+uW+dsyCkITIVvpXpA+R0q1NW
apeDUhE5qPe1W+mSxVN7U429kynPJP9Ce7K+3lvigucfIFYO8LnqIFmvIzPf9fiXEFyCLz9R0zCt
c3Ti9wVLQxFaXbnDGIy1qK1A9RXBhpkMSUlI29Br+Cm5Zv7dZF13IyqQuWIhZdN/I+B36S6PEtdd
w+tjuTSNa+g0LrorH6+oAAMXS3HZqpgNbL9eUW+41YA7c8OiZ0fLbM+K+oaW0+DIYwqmf+ipGvpq
85NxD27dwUmTAYwMRA61pF50DBjnFbr0wWwdPiNpCok/82MnBfYNqMFo43McRQkfFXdfZDPfsIN6
gY8FhFic6Xp00G6r38UVgEmAVu+WIID64fIznzAJd5SoQkdk3mWq6pNX6Gn0fnp7KTeC7oh2g3VJ
GAp8gAPsxjDH6HM275XRgFFL1yJ7JIzJ3mZ38NUiWSDNwKNmhHeLawjKpi1pouzF8ZIBHqyt4Y8r
0FE5J4bHYwHZVxfXMdHav+XL3VEY4C/VnpSVfPtunY2RUyVXS9eb1OwJE5yAQ4UmgXTktafzHDFK
Aij2hXpG1is8uSQerdjIsZbL+pt/xd3qAPemZpPxiKDMJmcsQJ67SKKD8s/fHt9uOPhgyWNDb5+2
LOS+dhBJxy8eMLfTQDFA+Jt7FyB/spGdbFY+o79CZAnxxrr9PYpJba0cy58bOi4fTTE1hbkcpgf8
4k4XpBmvN/VmwJXR95+Fo955iRjqcZzbLbz1N2wnmIylNMLSCo2Ou0v+H0aXLEYwJknpoqIGsA1E
qkpYtO6Ql0wFYn0jcNAbGFwVnM/GK8r6p1DJ1dzYaCMR3K6MQXfhQCrAcOPN7g1bJKnkMk92KBD/
WDHZAsN3nAV/btA3b3V3baeIB/g4DybxnjvYTQ6svrGxLzxGCM2ENyGy7PRyb4hYnJggUvSpACvg
GeAgDt3nEskfnJvEqwPGiIa0ze0N04z9+JcCgoFfL2icaUd2js8q+5LbMMKKDIxt2N4bG2qdGKIC
SzLDmM52caGVbiDBYhIN75iEFgPhni9YnSsYi/tVoYNUZOexYTH75K2QFU46rjCExv/7chA1oI0O
zXG0UofEbZ+FFpaGPCIQbiV/8Gf5zj9L25K2EhV0GalAFnrraDBtpkVt//o2L927xmxNlui0j3ib
dyb6qMvefkf0V/p5UqMCVlFktzBIIpxwVi1LUU8MLSQ3uPgvnWDgATdCogaMSw2SfPKxE1Hi2rzQ
Tv0rXjRpIuhH7Qoznam4JTfD90Kh5T0UtxFC/6O9SmfaYYaAlube2yKcsC3D46lrl8tCTWIf2DiS
Xv0z2SDu4aCILOqSwXn7mc2n2+jCo7Ohij36+M2JxYIGmvWc75L5y4a7ZskxDt+664ML8iNjEstK
RKyUYWI5JjETWbooqoQGtNnJCEyqaKgeeL3fkEgXmhKczU9WCpBcpOv3Zj2/vEMgoGFy7zTAu3Qc
CVSXKJo4mu3pIyKn4ALQoj1Uglp0HwioD4E9VNPPJowiyqy4JFAmI4YozcmQRj9Y0At/27dc23gE
7SasyB8wLrr6p37EwlPMOMWCu8goI5fN241yFuxFZKS309Rl92vwxJ2XpkVHK1kLq8HXVBjn8pwu
zTNf5D+W2ZxG4fsDj1tsQMOVn84HF0J3FmyCx9HHcWQ+4cIvXbvln75rMinHaWfzI+cgPCLdO+IX
pLxaLxqNLzxF7VAw/Gd5HyLvCzlGBsAZwzaSE3Z0ap6jiQGeKUZRMcoUTRu5N3C3z8H8zK31LIdf
eVnkbNKK30qahSmRyLjahW3RC5WuAUVCjIJ3ImoD5OE3XknpqkHT2GD8Rc7sBmD/9vo+bAQL+R92
fSPhMAWZ7p5unmrhTSJbi5PuZLHpziOzeEcfy7qQsJGH8qi+FtkkAWQcDCgJdAEt7STVoSDEAMmy
T3GFn29A4Ed6F7Vxw8dSD6bW7DZeUDlxbRCg+R9WUzqj/6SjyoJ1dsVo5ZObEJmff1w+NHXhWa7o
s0hFMopB5L3Zhy3blKfg0yBi4oKSIBh6up0uwzacxRVv93u3wHR3PoaAQjZoeHvAo+1zBUJnZCW4
8i71iRxAYGPaUEtxt+/r5NDI/osIZe//ujdljXqbTmmB4D/s9nOMbYkwY1Hyu9aYhCG457vx/vdX
B9RDXGF2oeIeRRVA7dqdEBKoMxE1PMUCNrn+yK123M/RTGlatEPNdGWJpphmngkbGBq9F6Gc/A/n
ukbRG8s33i5pJdOZtXS/Ep4ryJyiynZUPEOWMAAUyfgKPVcKz7wDhD7D7Lc+RbjPUiReDjE3evBK
WaBWlX50mAykfI4Yw7v58w717X8RRV3En3kQ/U0pQsDIVvj9/JYVqAMRmrtqjJk3soMZFFdBWlNZ
10U0oUVnlg0DefOUmnEUb627Lm/htFffCT8aZxOrogJsUMmtAUWsX6p7Rp9HbClVEZRB5hqeGek9
BUPp/tKpx74uvghGy7JBK9SSV30Hk99DPoB8FuoDav3EGYcm/ZEYFRzM8OocQ9tZqjxDIe+JjuPz
o6lQUBLh99Yz0tO70QkhrFKoiyyLX3Puft6lu2rxF2WgUTHCDg0WrUy3DgV1oFFO0EZQ+/RywTp+
43SwFF/X9yFcel5ZFOMZpW8zHkzQhpt3LGwGNzwT3edeaw+SSgQrHco8W4K88eIWWHsckNyA/5B/
XEk/aEcFrNu4s9M0ACWr5NsurujKnFpSVjb1KvGql3QT+5Qq7xCNczaX0FABfoYklB5Le7yHPi61
p7PtahTdTqp0SKTyenF3sSvWyRmFXN5ErCN7gxkVy26goxCrrJTZ6v66uU8CkkUBYI05Tjqj4L+w
6tnq9p7Kq4eMcnSy8SA7WcEJAwvB0Y6DmG4S8/QxMzOSA6TZcOBnm7tJIOldRCo+nPhXy7PyCiYe
3/cz/rcvHN8m+kRKKfqMyIg5kF1c5kSJ2F+trX2qafwrpYNxgqj/FHMQroXiIoFqMwF8CE+0K5ro
kCItMh2wZ4qUIjfttzjRB9H5dfl7jPgVWypkIxxQnvsmyXBY+1UHKr1QxxPyV/y9Fgd52hprI99d
erQ40PNJSSiqcMz4nX7Frt6Ts3QDKvcZ/aaxLMafBxZUvBa2xBK2SV+RnN2Bop0F5NSDt8B5FG6N
nF9NmR/S1KDS6QYTsoOJHPyM8blDmgjiIFH/N12OXGaBgbAZueiocDM/I6YVaI0FW65/+TyJPCTc
w+DM+3iwP0pcDEdPVZBmGun3njEGXY1kn13hh2nyj8CODADW7F+KZbZ5eu/HkU3FOD2IGF6yAc52
y4v415InITBlwO/LadhadKxYwHO+CSJBRslrSx3zF+EhobfMFdgtGpPoPm/sV6tE+/Ov+3RRl5wK
UWP04HS21HMpLlsjeKQTqqdzu7/KglyJ/Am8h3PafuUX4Q9wCQ1XaEp2S+9UJKjDRibLD9K8eSG8
/g3naJ6zYodkVznehi+YSmFy5UOB6hjDzU2QR0cmjnyIcN8Ai/VoexreECdRTHXsSd4g8+UhYeX3
NWtaHc5BN703PTHpSwgU7IpsAfTKhIcuk/w5cR0iOaYvEkbP64f4UnwOPQHp2h3ezHENivmVbOex
9Toqws95IMbEXez1d55vNBS0E2EbHF/2VodEqY5o6wJ8bhghsA/jSu9ZWNtKGyLrHx8OCMmuQ9tD
4fdGDK7TBE4+GJOjaf6n3kjWa29q5rIbRMYE5WDCx8MdHGjKi5WXqgvrD8rJnLkxhphxr09hKM5D
B2VJFc0SXptJFQisaKwCNcH8/NqwT07QWvQXXhmt3Xq5kQGhyKv64mvbhyD0jOzj9tAUrnRMqq/i
cJnIuc+04FT30BHnFjK0x9h1qgPUJv/k2jU48hqFj+P18UjkUGn0GW+FY+bFeIxXYrGHESBNzZmI
Qo0Qk5xVvp3+3reIExzfY3iCFXusZAwnJcYqqPTbA0PXwSMKfR6/Hd3xGLtqZ9D55VG+RdBBEopq
OJzUmLrE8fQxafaeAGLZGwXyBu9cOh6Zuw5oAEedtdRsPQEdd7mpyn3/XaJTGIyQ2RmJrp1XpNMy
kAflvfG9afOzDNJJBnpG4Glz0Xi5Me0jUyEigz5oIBPz/9Z8lBD1QUvH8EXUdHBaRGmMjZ047MZF
r3kZTtOL7YeWlUkWk8GON88yttGptEws86AQnK0nbncM74V4cTW37nDe3gBY03apJQ+1+FLCHtcI
eE5Maly+/BksYCjGefELpj7uPqCt4WTNnoDatsXICZ2TjuYQisSju77QfNiRTaz0HNh+45MUkAWJ
Bt+mfkEodsqyo1RA//5PguNyBQdpyMPRkGXFFuT0rNQxfoQsnWkW7WMGZDoTav4pHfL7iVJo71Fn
nXS7LXG5giRk/dvCjxYmRhceH7ZQ3CBfGaBNwOSmV1b/qpSBgtxwGRHkmrAS2gnYL1imaYOe2EAk
7qcQq6wXwpmWab3EQBC1GGHAaikI4z8UxPdcpEhcGFnRwNE5MbPSgR3+TznCcwkTMKqUkDhDkOeu
YkwjJ09wdtT1667je0paofGinWVA+I3cC+7tfCS0GLLQNd/IrRf2/c9PyTO4XoUYefEQWdaMyd4S
Ri25rv5Ul/tOCJp86s/4y1MZA6gZEm0RjlhIiX0As0dNvrhmgyDzW7HgzPYHRyulrrvxPpFcQK0t
usCEG25m3FoSdDACZbFVAiG1tbx5bomcQn2suVTjydtORuSxPtQADCjsugD3c4u5EI5FktcmR7LZ
zOeQsBH6mJ9hLCy6QXYbsmysYbndC5MJvUqGinlRqvRxaIolJKM4kXIP5OAfaV3miQncdZ79OOqo
zkawhVufx+CWYVaSfSUWgdUuwfkux3T7dU+I7CUEzz6T5hMAyuFhH3PtN1W8CrvtNg2BdpbZJYeL
KEy1zoUg3DNX3LVu5aIuU+5SCtDeB15G4HfD7rZJdrMdE5gZSPmlDhkdLrJYzl/glUMD4PIXoQIN
EP/Swt2IKgX8weoeZFCkBHD6KNiMWkb+SD64RFznNsqZ2pIYyZvMJ+OzURqt+0liGfJAZXHEddG4
UNJntl4e3qrBCHbE9ekYiAiAao/JW/d0PkCYHqm+WeB2Qp/v8AgtZFQ0uH/HjcUqOoiPunYA7Ra+
ELVZQV6k8PuHApen/eVPpsn6h2Z4A8fJ0EaJGGdrrHxvj6OzinrPqrrBFZEPj0LaX2jQzpWwhGiq
U1kKeMpzJsEdDC4cTngjjdmZKqoLRM6vWGavabtvNh/cRVhXI+PgvuN1N4KqOFXeIiUGm/CVLj3T
5OLNq17kzB7FHmSzFOwCh3LZIkzdEDjlzg0ks6w2SBFa/2JkVQ3lAUKIX5xmYWJv6PRwJRnYzC6i
Zbou0BW9Jh6Vf+H54Ya5+rLHVQwxPO0CB62HGNYdubG0TjV/My29YhafFYYIg5wnYfMWnR/OA9Gt
84XwbV8zfqh1/uV62KZuzFVSuV17ZpZUHNR7LByFXSQUCjKxbmT2BYyfgBTXjkkH/u/02gPqrl0D
8vMTYfslkgnqbGJ/BgZYNgb+y31OvlXPUMdiQAB4tN4wLs9iWJyhyGUaUjSk5JGJUxiNy52Txvbp
l6VQ779EB4pMtLjlZl77x0DGQgHgLwPrQxRUOEMy0DA4s2Xid4dNxQd7K5gcSudVwm4TJ3YcObMb
jj8nYPhTqc4pMXu0QhSN5/PfFclqTSIGZV380CctHq/Wp1J1VLtEfulXQrtt/vmEhNSpaXxIyGHE
f8OuMaOqSWRDRdCCA+HZ0axjV645d98fBfzOi/UGtmDj8c8GlgJhJ8Y/A1A8pMHxgsGnItC8/xpi
ts3gFDwpacWtJRFkjQ70FB1ZQjIkevkYPhcG/FEYUEykOz9M6mQ2b3ma6u5pUZQuH5AB/fPAvFb/
3Wu8LwE8dl5vHMAbn3vwgZwL9SuFpI1d3SKTtDmdw0MSMnqX6+9bUFfFTGjR7kDXb56wg+HNf19o
+t/oCEz5wmYhGZyTrkhZL8vaD3qPBTs9nmU+SGmaW9XPByYHpMhmWsnyiV0MAK1p17munJgaWf0Z
mZR+AEr5h+lW/DmCimnyohAXtPxOt5BTMfPQ+Wi+bp88O9f5163FzLjBXKmJ8Sh3LG0RbRzxxdvv
4wGV4Q/3f7+L8qKc80zjijghBUuG201ReIfPwZBDlPAJYbcoprQ9mHJhgZDl5YFNxCp78q1MJt0t
ZzUBDcO8sHPK4g9f5o4EIO6hHICksiWJfMJKWN1ZMNmh6O3C03K5TMsnEAENw/sp8gmBXFB3C9ZB
VICWJwDQRoq2bbCbdMbk4i/uSjbmJuB07fjd6ZTHx3ycbqpQnUmZ+VDYvPMWWJR/8MGNC/X0gklQ
UrXzyn4YSIqcqFC416Qv5SaD8rqLLx76E0ARSfrLRe5KtJf3XxR4DMsz3uIJWm9zf/JY9MEgDrCz
00Qo4qizGy5FtsIEYJa245/N7g9dmkcG4qln7dFbEiVfsnyaz0B3xsxICrX88Owz8XN4vXVEWqHq
zcyqBiq6wbr6ziVbFBBfDEket9lpp/CAi6UimgZj9ZwmywQiB5XD3UKXREYQ8Z4/7NPAzftJg8TS
S9UcAxyku7m3eYvurogqtYVo/oYROyB925+ICb0gqRnfxAgzKVbR8TZ914RD90quviNM4vo2NM3W
mKR1EZHDgdAyOMW5iuOtFv3mTZTIkvqTeelv+TphCRRZSWEnIquONWkTjSowhN6EQNoCuacQvxCD
dcVFdnsVgpvp9ieolly7FOJ9NwgkZGpBGOKvKRMe+IEDFmW+Y6/u2l96KDtr1j4ziYE++pdCsWAm
T7R401ENLxoj2Uk8Huc9Zjg+bI9PXP2RKqIB354Y8XvKsPERzPt1KLxk/AxU1eRQMIwzBPd5G0In
DAUcvawn+kyCSNLDRSPoI7aWrKGpACgnOqBPwD55UQZFrEOiDGo/mI3Z8375r0CRacgXE1r70h3b
9w2RZTgjUAkD0ixh8ZQCBudORqV4rE03ZmHGt7tOLh2ridWDQyxOnQQHraikIXUbgLgUn5dvi3QK
PEuCh8oBghl8X0MOPv+BUn4jtl2b2hODf2plTBTOxX8rRy6u5TXlyQG9NekP3I5Xlbrgw4LksAtz
F7j8XRCYtzkyxenbq6p+VE3dJlsNs4KCXEyNOeiJSxfJKiqeW9lZowl2UMGHoeKWBIa8rl4nmjDi
makJDq2fLC6qMMPZPcp/54hfZ5X0ynhPsPkhMsfodtlAa5De4EhR1EMPMZ3e7k2otQ8MBgVE163K
NsszrQwzqGe7S0o/emKC4Ql9/LJM48TcY111o41foicFS74HMoljmEwtP+jXZ4hY2TvMFgaQaHwf
4qFAdnyj1NjjDUqSHOO4zXqRo7JVt9DW5dByCSJqYU7mV+MXo/U+pmZuHRj6k/ZsYSv+RBajvB7A
/kkYi85ym5C//tphQvS0viJhDC0MlW0i4Z+8n1YIcueXarZLqtubK1/ivtSSLftPXHtI5VQZknWD
q4kA4c8hN4ofsXkiq574iGCn7iCj9SJMhIZZNTnuGWXmm9MXvUlrh0Cj+7F7hYL1SKLg0XK29V3N
K/z1WgmW2iyYJuuD4kYlgxYkP48ppARCcwPe2orsxuq6E6pUeJwcsEDoAdNnMjCfzlJY5PfPaSeU
vnI1KPDdxargVJ3kKV6pMEVwyaUXHpvCioiovBmcEq63Ku9EJK4DKGy9RAm5sEp52Kf6JdnfC9av
/SLaeS/u95ZQkqaCU0uHqEOTLh4klNvGMCiQyCAGhMYhRXVLFqiJN5Dq5Gzm4DlZC4V9xwsvSNbE
4M2zXotUHe//g6xqYdTV2U8iG3Mgz06j+6K2NnfB20O2FKwgltP59iqITGA7cnl28P4DpztD7swF
nF8ufXPhmta2T+9PAJPeNnsbu94rYfc+1rukabLUthfVqCK/8QoLzexaYVxZONil0b6RlqfGYJJc
Lz3Zc6FqbMJfkDAe3Mhf3sNlEc/aHkCRJldsYAqE+OnMLY4L30PhFL2O3ro/mbHjOlvjs9BvlY5b
5GC3sj2ANWn2ULK8t3kUAZUjKU7HGVABWg18goSyB2thN+yZcpRuh6a6pHLom9mq5ROrU7K8OxHe
vHij9nVHDK8mNSnyrYdPshloNzKxl/9JDCKDQF0gv9wZj/O6G6qd0AUFnaZYUx8OWjIVM+CYhpyV
SYCmniDxm+XynpMsJ6FAXLAu4Wht20t1xNzakw8BV6GiyQIzhe3UlMJVPymez9cU6PELucM09/DH
gEXzkRKrAwX7e3kRYDFQCUYxy+oopU6N9VX7o1zRWYn8YSSuZtiEu2Z03mxqf6ml5wWQmsbThKg0
a1pMRD4nwlU7aaa8QbwE5O/PywOFpBwLc2aDolyp/p/WIJpmJXwmpfrI/YjOmD+7+RkFjxZCKybS
saOYYqF6XKAwJ4fQFVgVtBAJ5xLjDee/DI7yikr2P1961tSc0yIFnwrL4XOttlb1G5GvpqV7shQg
VD+YTGX6nPKqihmWZQACIaJiyXp0l9/WfH7TrW6ilPe+sa5l9mz5J5sqsWT37Zobfa8iaR0KjINb
NSfbFktZw6EkvvHrrVlnjxG6bi65K5aVUGb39iOEViAPxuLWZMXOQ6lMfd39N+qtQbzD5BG74xZI
W1dn+aV15x+iC28XipRhxIujSR2SA/8MbrNW0gTrjSqb9TtDzUx6CsxgekDM1w0fi0BPTQ11zsPT
QZASOkwDdiAdrtUrf5G7jYjzwI5Aw+lYrdqBbODMOj2mKUeFfVX37cwzyHqdr0u60npj44lKHYAG
KcWUna9myYAVoPDfYT3/irXu/zoXnwb0SMvSGxQVqzutf0AYt8URg99CqPnpUQTFgnR4UqcAIQ3z
z6xm8xoeLk1Z8XXYtGmLFUOC71UyAVuIVMJGxGG3kUlSfTvZSJl+KqZriMo8tKFXMMFxQllKZ+F3
Lysi8OFagE+P+k3FKhuSwta6Fu0EfhLNm/0njoxwg8ZJ6lMkLmpkyxiwrIDAVq4uPJeiNnazkbgV
ULoxcisF7G+tYphhw0QuV97oruW+MKQQEr387bH+n1FVMF5cwW4mXgbMoU8MJS0nf2YFV/rW3csd
I4bG8AhhA+62kFdJnZG/LGDH2T+REu4ldDIeZpyKscUeQ4tlnklrNLtYdl03NXz//HXFXo7gNCwf
h7MpU8foWXf/xMe1AxSO6zuPtEsBMipjnU2mBnbz8iUCI18xmdsYvyJwVCOT9DcDoN4520a1QgdQ
Kw/N2ci9TcehN3Kxl8sly+HsG8M/55pu0QzTqdyKDim7MSUiIBv59R/NHC7J1zPsgqTbR0gSt8SH
T5EvCVXfNe2ip016yCzDmmAf0Tc2f45bD4diGgZRvNw0I2+2OYG6TtVZufC9GR/21YqiYoNfNd9H
bRBe2NQ31ZqC7n9C082SVWaipIC6kHMFUseMn/pXWVTojYAnHkwJL+po3A2uyQUi65MsO5suaVvO
jgA0Y3sN6cILNpZ6yMDQPIOpAnpzWOiM1x8jig7paIf5wLjwbAUmJvGvZtBt1H+CYLbeqO2QyY4D
QZSiLIrf0SiurlPzZomy1/MIoX/OgcahcXXyejiPyOoYPShShZnvl2aZTukHC4NRwRQPhb7PipnW
TBLS4jxcxCx8OfZgZd9WUeegs5S/Udgxidl63KxMEVPnENgqhrNdV6KtmdFZb3ZLlhgJDfEeNZOv
A8ghj15GLW0DeO0zIVu7XThMjVi4HiwCTi4v1/awYbPliNWsTLy8etmkU4p3BhyuaXx7vmsniiGA
34EwTFCDJ62oJUevbR+4kIcXTpFyUQ+wGub8UUOs4GrjBDK55h/7dy5gSTG2Di8Ec2YBBFwxtGja
SKbRW+OHX8cOW7P49duPa+V50RiaRzJnvL11D/SKwWhjwbaXL4c3dChIXBKMPvQsotIdM9stkjtb
frZKNdRM0DftDvJ2zdvx11z6Ueyq30GnuSbm2Wcrhu23kC9ZAlycUlEk6Ekby+R0ICeCJLLL3sS7
tbW1NLRIhzcuzjmtKa1Euu9qNw90pP+e0584UFuq61gmAo0fysIWsjWDe+xTtwTwUGO1LhUTzKfD
lDiUwMEPtRuf0lslVFIdftuqc+y2HmzIZphpjyLQ42kXexUTup8MtxBr15WQCjta/8eqnPTn7SKz
em1rck2np/4he9cG9qacxcpqNnNMBSJrQaQUp8P3Igkxv2YptXppaJlP9yvbeRN3XPP7jG7Z0lh4
rLMoncx0pGBNpR4c2epnpTYs7SeRLVODLPFq6dfKhaASVuhfYKxevAE/qruO/lXFQA4QjpITpQaP
89/lWUmPYIkFzF+vEJKqBW6/o44POt6uxqn2BFfwsaoBPh4pjIg5otZESC9G7RbMXEVK+fSASulT
nRpALAZ+yhpDtlVwRdpcGG+zdmdjyVqknxBo+4IlDg1AQX0Y+e8Wb6m4HH8G7klQTcsawqVPXx5B
MUCkzJyKFvbr8MT1Au8Rep0ohxpZVyhXjJk9/wnEywqdDlS/BZjDiQQ0BkXqBNKKAT+jwUtUYq34
vvaheVENa5emXHVVIfQNr3wug2Sk/TM4XPORYgDKUlptVL03qyQOM/fQoxv9l46an1JXncG/fTn9
B9ib5RNQI5iFgIFSMES4h1/mqXxZ91Xy1ptWv8rgL+Y6X8+V6HzpgDPcZWTBnWNam9crSAYeWkZG
BBhegCN5M4td4VterAO2l8hrrMk7TFX2BbCWy5qBJbhdo5phbUIJ2UqDMYdg7M3XByPvXnU7cOxM
ez04eLNsQAm1tBR9BERjFxsq6zuJjFZvbtAL1CJE4302Wc+RSc0eZu/zqfIO95T7mInNnizkQhDt
9vn9uiP19nSCpnc8kH9dNcWV9edy9x/xTpQTKSazVKYHhZArDvyvfDhnOo/v7rB61FrFsBfEJSkz
yXwzdc1X+c9YBvCHZMB2yr8DP5g84gUT78nw4bDhpkIG/v1x3827bl4Jbp7EWUMT1RblryUvvlNa
RREB3Ppt4cWJQf4j3AqYXs4c7Jo6xzhAVH/vfaHiXGn5MKqTR8WntJPCfB6H2JQHAH62wPVVtbeL
xJznzuZrjWSjSKid9gmJ4B5tRdrlll7jtWrqZ6YeMTB69vHdXKkyPOS1IzVbkbvPYMI4WPKKkJTH
duuMYNq7hz7JI6d2WePzUBXpExbAf71cafgvBzPQ5D7vgYZCjJ+QjzRxH+o9Qa0SlEXKdA6F620x
hn4WyuDBcOjZg4WXvOtjdCO9L+mfcmHU1cmLJEdaP8rTIHUeGoGTWNqZxlJqDQT9zsNiqrv/ZnPS
g0A5WcJhFxqj0PT52mnQ53ryP8qS3TYV7zEcmdJ+O4tlg/XApWAGfbD/yEtvVZZHP7dQT0p2MW7i
PBCanelt+oKiyXTHWvT+JfXrwMdQP3XLrnoxMkWwVBq0okXIeh6bo6HecXMwAZeIDca783YPIpXk
xK8N7qaUYtZcAPiEX3vpur5bPOno8VR552HOf5DuTyyDEcLqbMkEzE3OVqA6G/00mHf/vFKvGAjH
Eyvzp1TiW8mgo4J5jCUBLD89/CXGUjM9l8jhSGurrEWtdeg3O+d0hRI/BxRioJ2R7BbOXBqPn0gY
Kzrn2wpQD/zmver3tnaDU2436EVnKAPtSFhg4jY/hKMSA3C7TKDeYXFiWaLWkAJkFZCcUk8jjZAy
9t71DzVbCHpWB2+W5JWHyNZIZqdSV3u6Ai7ImabV39I0o3uXRFPg4zKwQSiNSmgwNsB8HxtLglV3
wB5ikkjcfC6+3grIKdZIPR3dJU/W2caRX9lpsw+7X6epvXiCwvHgAwEBO44b4zEvS4LeuNLDJ0yM
yZbmBoT3ezZ1Y5RU4gMSRFZ4f+mM6t9t1dEy//C6tBAe1gnynwduafO/RVJ18G3UxFOwEvVkZRv7
aDrhVZ7LGzu8/ALjzh3tXcVhTcVfl55UW79XwSFETjHQYX8wyr4Lo15jZClQi8fGhWrU2jSKK9ee
VSmS784XMRIdepH9NtyxyvVW8q7r7+bG4J5vChBEdvb51R8vZoGc3In5RSk/t5GOiqJkbqBUb8St
8sfUA1VVLxfAKZuxKQhvi1dKQDcFh8gLaYUnH0Kh38kJEFH3BKs673epOEzkRWUasy1dbdFBl5oF
V/csSrunZmhnDe0A1kRFXWlWBRr5WbIdQAh7wOUyusId0MekU9C6mveQCxY/aWjedvNTQzhyt+rP
LdPA9Mdid07RSNLqWpAxH3ybZskiCwN87Bmm56X/GdG5AvotCfu88Ap19FT9gqO2KOBLh9Ef7pc3
zTuPyMM3k9NBecKPVHzLL0vlow8iQzL+HdSBO3Z4qTne+tMzVExvZamuJLIvd9OZLjYZpNtvmWv9
UjZ7QuUJz9S2JzluJE1dLo66vJVixUeZU1eFuKN5ZOQ0w5dSgKBz8GLj5LjTW2+FTdDNgLI2pUwg
hFZDPaILXaJJXtl4X7lRZaPAX0xdZVLcNEAsS8cdU3txFctS16tlqDsHSHHw9awTuhonDJKTXzPq
UczA7pL9ryTdg45WgnrxmRaovR3yt/CBj25fW5K2BQYEmxYxk9VGUuVYH5al13jdnlFHFQlNfKYU
RQgbckRXZRUPinPTkGjl//XG8a7Ystl4H9WSPcvXaIheKYGrEUfFSno8n8U7hJmmcL5GgKDXV8RS
kr1Ui6AEByb+QprqbtOSP2HP0jhweUmeNmrGd7FvNzyfSMVbXtu7BOn5Osjw0aTptB3WdGaBxq7R
+KwBXBmd+Tro9KMBxQXZJG2UwpVKomx0I4X7sEu/vHES+XDPbJXJYPSPUrjmuqs/fOLqJZCkeD4F
fGfFYoFo+3dfHbujj6ssTvVmBnR15Y7D9dW80fMPGYickfYWO7S9udW7Zj7ntv9ScZFLR7VQiaL/
1wdTu+4WTaaDsoxjs2Dz8AwzW7BO1Bjb+MRU/2CAIuZuR6gM1AM3rNKu7deyZCPVC6xWPArU0P1X
kBQAz+aIRzKDnfZ1x081g2d0wvAcHEZK5alj7qG3JZ45Wj++ziruHgYSt+2Hra6OdXykKM8IyEDp
BLu3vKLyniKDqnxsxZNliDq13DCC0na8DUG7plblCMqTBznsf+helXW3d4MiWE8mliThVIVFf166
LPE5YrhvNGYldgZWIiwFZ1sncS2FPMJB//L5vXHm85O8xRTkM5eCzmNGSN0D2YytJH4SyHz0Wt2p
CnvDF9MP9EJCGQU2fIIa/zztz2S4DGxQD8gop/LndWBYVSFWAG03MfE1+FxPVbr/cGOwPYQ1Sv4G
6en2WX8NPLijJOFt8z2xQjFUIb0vOsG5p+Th6wYEKcAgWv5AipQfrOf+HCVny0xpnCn9VIN2b3Wj
P62j+bFW28X7GRLM5VAQNdBVYwdmJQiHT9CClveLdyrzB84S2DMd3TMHx4wvKLWZvyUHeb8spHJm
VlURmMDAbR8GDRqBnwVfuOaFmI/sapjDtPKKqtti0WpfQMILGUbcf6he2QQWXOX/KmxkjaXcGpCc
Q5bBl9r/KnOTQr2l0JFChKJlMKukcZxSxwbU7bcbyWWu7KyoFx/1TrjBjpo4ejqy0hrqRaA4ExP4
9kLYv5ofK+KLdvmMio5GsL78lhfXI4ZQTM9S+WQxchDcTJb8BvqhAr9YoP3YwRHjfeCwXU7sp32H
HQWVafNuycLkmC5EpX794uFcFHxhGUbSt++nzQ31+JKl9Z+utgoHvhxEoMeb8U5Wsp8rGGaTafA0
Ri58ngTBJnhAEJ58pBhSS6u75K/phMv7wAlUdvdQWneNdorzSZGeb5YpNn51M2hwtITL7GtFdCqH
4wgV+avkqxhpsYR19e/h0eWWrkC2yjmn3G0YIlrh6VYGRUL8j3e/1UX+3YW2Gmf4bqJqtnkxo1Fz
L5El1fmRL2iaOQOs2SmNvt+i3uSHBzFw1hNH85nWsYPv4R2hW/zyOZLq6A3Z2j830a9uDL+Zbp90
g+MMrzNODwvgA5ggzsXsC7y1VvvwX440q9idTGEpZty+qZsC4Brfdmyf+fFBh63tLDJ2yItpZF8N
f51jAge5ZcjvhsjMTCaCaleaJn67NmqvM4gSk27DmDxBtl18wWaYLz4JIMsABMLeTJdBZmnHn4fE
rS3zpFsiOO5EQfLNI6HUdWVx3NxNpN0K7xpYxyiPvOXZQgsCGhju4Zvhztrimoj5EhceoygB7spF
XplGGs2UhgEDiUdk9r3RgqGQCGYNYoT16JX2yxMkCGtuPnk1iGf1PIfdriGZ9mbcT/uHpFoMN4Kx
c7s5mIQoDfVYyYRNx5sMlxmcjwV1lRmZj0oukSGVh39MI/GbTqp1VBEC2o7FSVzlmVQ94QaUH1UP
8R3KJT6L8/TZ6foEr031VZ4rMEnnbdusGKyfkj4iN5TXb+ImjRsfXm+TJoBxTMVjS5ewHzR6FW56
TW04t0K5iJ8QxoV3TIH7nLk6OkYWUX9U2idr+LF7eldbk8uT5twwYtQC/92+wLliKMDQvFUv88Wr
7k/iEYfLu9B25ww1xMgncg+CXHr+YSOZgJkpMoE3Bj5oRNUJkF9URXV5tHY2FQkbySBtpKIh9/Ef
FT8jzg3BMCQZOr7O0r9zmleOV4BNsfM/41UqLViSVZlTjTwuStGum+UWZWiQuwjAdxEYvPytDhfN
DY3C8d8iSLkJtqoXuKzaVPPG+96rr7fzZo3h5NEuv/TPlkenBzf3mvM+C1i+szw7/lYqVeGyAlCl
siE9N4jUMDVQQG/NyEz3n68n1ot6hlS6M8H3cPB2a6r32RW/Iycr2f40hTVwMDuLj4ydSHdM3jI1
uAkxSUUvJ3AF4Po6I5taBbFyDPhAB4E1RG9MGweMSi43P8VvHYHs//lu9tUT6uTiyrpX9AX/Hbsk
bJFTT3/84FsbN2QRhzysEAUmbXuXWpd9GmKJcpE+i9iKSfvf8pi6ZTNpE2kdkaCMLPfKDl0pvzKm
sBcwg4nPvX8IfLuo2rsDWj7eCgPl9tq3xOeZh7x0KkZCaxfuiZZlAH4a6hQ7GbELc59amut+S2WD
hsVf8DqBUkl7gfaT+t40aZy9G4PckPnFIc7X8FK+JFL40lmt2WSyN5GCtAKO4QVh/9U7JZ0po+Tp
2qQmRES1zBTdmvM+NELgysVzabexXmgvKdQq6c/blQ/jS1PeIkfZxz2sOKWeOuNXox3bwFDVL5vN
QQNWfJHVYFVxSAk3JZeAyWpVEFIDkTo12yQBrDCRHd0XlKHm8r9k3ccVN8gSfKvBj+P8A4wOqre6
Fe4VMnCd1iuG4Caa+LUiv1i+FX2vREbnaLaarOuQY6MSbsHXqNoppbmeV3rhyu2fZQz146FCmymS
Jo1KXzjyruaQGiEeXHRnKQdiQKyOm5T5we2438lLa8nHs6p8Z5D81dDqir0tivxzzC2tAeoOgZMD
uo3ucH242DbS5IviDenbOU17A/U3ECuu+4uWl6CsRa3ipXTyb16NLxcrlXMUdXcPz4HWAAur0YWv
uh77b4NGQUG9VXjh36Hio/LVrkv/XeoqqWWXXMDdMXlX8ry8uu9fczyfwBi9asrlTHiJ9AsyD+zH
7F+UR4qflNh4Pbx9zD2YRupet+OzAVhEHyVGwSiaLkO/C1Jkg7iglR6dZpmBxqOlotVGML1Sw93K
CY2Unk4nKKput55HbN2l5TWBsybJGlvwtZrMmbXIkHI1C0Oiqmr+XevTqDXb/bku59yiWg9W57rM
3pxqqAxCPkmPdyUDe/pY9JMWp3q//ed1uWUqI7IOK5jBAEpKIhMDLNe9h8H1ePZh7kPf6rKe0fHY
ag33wZfu4b2w09QWt+vHSevcv66LP8/m0J5KWZICjxclCChsxeDHjxtsSfywor4sJTK8iR/zWs/o
cdUr+2msTULDTz9knw1TUrCHlPQwXu0PKOZfpv+GuLu5dGwETM05XpuP2ZW94WsR9a/NOqRr/N8S
TVysj9/6+N3F9MDz8iLrEJb94o/lPob1FvSJqGt8YFYAdcfdmhgBMgs9FACdKhkwIiQcdt4Vw/Fl
w+U4rPM2XiwsfxVHTupe8o5LOIcfTjtqrhgDFqyIn2dkysytJliTPtWmhjKg5JZXvGcSn1dJqJfz
0Zo81FpGpcoAj1l+tRZQd5MoubNMRKsqiQxl6vRiBYqN3Wmq8wog8ZpflPx/BxmNBNUi4JIxrs6y
vdI5wVJiz3Je54yj7C7p5Sr4hUdtBV3BYoOXVuKSMwPCbD/BkcXhSK1+ug2Sltn59PZ3x22LJ3zo
qwackpb8cGGx+OQ+s/Cih9b9Es9kTToBcoCQo8uDXrrgBGZr4JRYtH2qrvBW40tK6yD58br/RR7B
L5GEJXEhmDyrW/Rv8lMBZX9EC4oC5yUQzaiQfvk3psvOo4+VhTfFSsvYwe1fB85ttraHpO3u/CEL
bW77WzlpnCQz/e1vjUf1j/hC0e1ydNg3HQLQDcyivOOPmQSTpNqf9RlFNStEb8CcG4IJLaQEI1Lb
FdBFnM279I2lg9HUIlSTZxqjR2DdgOGFOlacthPRagN8Drf62u4dbgbUb1+B1dZc8apgAPXt1Gq9
cC6b3WwlN4uVkt5gKb3EZCAHiTykwL3wK3MDSN6s4dqgF39WJuPoV0eGgfSrsDiEp+cnO5CaqqfS
2Sg9hEXBo3G7GcxmiJRb365Y1ImzjG5wn+GsJh0SNWl99sUpV4UN2HHac945qhkh6IV30vs3y1DG
cZpskWp66+EM7ZxM01HPGH37F3jKdwS1l+nPHx6mnHTzORLch3jGaLnwe+CKNHmAT245kNXiIYrE
3aDTPOMhHjsVok5OGbKroYVwDf3o5KL4FrOcD9BVjTA926UZnB8uZAOT9jtK2yJBURQ+n6FmErWQ
mc7maj5FL0WnoqCHX2rUgwvVOougV+E9Vn330SaPCrsi7r83zdZPIkB6V0HvzFzXCbl9wHjvTS86
w5l5tfPKcL83/WZba5vGgT65rVkZ1C+B2kehxyKUgCMwpLwnDuhWtSsCA7B2KGnKzl2/z9gH+xZz
DFZ8HcFiCaKdQ65DBbd6+cKUphAai2iEoE+WhUuXtvcZrUNH+dIgLD7RA0ktR1eegllnNUwtaqxe
XC7NR0NQDyIL+f67du9Ma09mIW5uCv+xXpmXD9vGIs2MpZE1U/z7ihSW0HTaY4gbb+W8XN8QLbeT
9sBFBv+mLamG0vvlySTZCiXglY+rddPwofizv5FSHeft5gQBi9FHPIJpsIQrrx70sEaVV+LFHiT9
e1LaRObHxlcRBAng+1LjMGUHD07h9ienb5VzNclHZiRsSqaAbDVXLROxr0ob5w6KBf11oKztvdr/
MAFbKh2u8zsg9YhvDlhKh8YRu/JEY/jhK8vR5xen3sJOUhe1GFo2pB8cBOmNVM1LUMKRWNRD2eTc
8TjYLv5XfxWMjXColklGwk1aEi/GgIe6QDDPVBuJ7Gxh5m/xJCH4wL+CWNuHBuDuJ7aagp8PqIoR
1dT+kHyh1kqWvSRDoKxRwfcoxi48bviU4Kdmt8jH/ZmG2LRE+UA/Or/U/pUfeuBggp16MEVa8cOs
PjMD7ES4L/gq5Gzivt5gvqr/kNQDUtiSsSoi+bRxDHds7UXbQczjtVJHh3/cwEI7eCBNpH3uWZ8U
wLgYdJAh49xfvnVAlIBuaPQTAK841pwoM6VvhSqlP2vQNcewYgu4EJkc35T3BwiwVeBmKU9lX5VU
iR9EtX97S/pndG+Gb6AwmZQXDyYvZ5SQ7H+tm/LfQIGS4xfUo8uGeDv5NR0PWmSnMCHHoT/BTF3S
+yg8uqb4A6F7QyWFVD21YXGxBQTeXw9ftzwkqOfAuSdj3jq5xvKeV+2DQ3Yvxqv5k+QLi3bUtWm5
f3yXmwQH+EtyWw8KGgjixl/1lbHiiQxJsiqN+2Tnx9aTalp+qC/cG+g0GquXJb38/HXu9NLBKXap
gEXX8ZMzqU6yH4bbRC3+u2SJjUV8iz9B+IAuYb1pKW+tgZzh3AHfZuvmkqZY3BPUeudZXhNtjGNs
ek0Bb6DXR8Vhimqi5qSA1ThDOj5ViuZ9I/T0VjoZtc9rO6Mvh7sUbnqb0LOcFR0gG/ovcVoobcPa
t3OJSjqUVgoR57aaUy9hyLU2s0ZdNab6S+/aonFjs6qWcDu5RVNkK3OYddIDBucVfcWjZbrpIvyr
HLWnLJVwUZvxiQylPvaB3gyE2KyDs5S352fzzqrI0iNOjrx5ruq1rw/5fPsVMNezyFV/V4xsjiV6
zo65Ca22OiHaFUG8S6xSTJhX6lrkUt81NOvyNeZMcIvf0m6bS+GOxk36kr0LlEOMbBv+kRa4gT4N
6CZeJ4jdV4HzVh5f0f++8RBeMx7ydp82+l7pP25herJSm3bFEqeNUTuE8Q0y/1YFmt7MuQFRVhtC
7yM9oZieRYPixuZ8yXh7x93u8fnvFFbY3q9YE02wIFCIRucX08uKMpGg95drpjACntaBcFWuAQi1
E7HDsRGVG8AUztMetMHU1+IsBXYzbkEJuR6Rm8q2E97RDOYRgip32u6/84DNS8hR2vx6XWUikTgd
cZE68ECazKKpJfKSw2uqXDREueQn9bjXsfmSweGMOym5SMdKVh5bp2R1cgxIJUVgEAUCSOh0PFZr
ovOcMZkCvgoEzmfAPLV81n7nAJHONFjvhGScKdXYklUxfCmp+nY5nPnV0j5n3V6VxJL/GwrGRV9Q
eFK9TRThgU/54rGTqKqDToq9kvMoVNtxP9noA5clMaZSxcOEMtU7n14Oym9W4q91wANqW6Uruk1f
3f9W4TrQta6ktqjInUK+GZqG5SKbfxp4mYX+HoQcQJ4O+7CP0VMjHarL2uMF862RshRlD/Mdb2Tq
a/EEUGK1e641vRuCtJ9GUEerv5tUAQtgoKwn/wWxYPKiuBmI93h22UJw7pA/JX8thfkTiZILwe/6
s7hxBBy0fkZDBk0n8mj+5ADkpwFeT5G9pcI/EKSvTzeZMCKosDVA/SmJqOdiOmsDawM87VEue5tZ
G+sIXvxZhDhmrJ/SSNnM/VNQXF1+8rGGGd+xWFmgm0HTb6HcrmiJziRUZNT1APl09HVME+Yv+UIF
AWf+W0U9/evCIm9baDhKcsNWW0DIsNf8kakDrB+h1Vik7oIOA6vYTY4ZeNVcogrECIlnRyi3b2OW
AdUh6ehDs792yCv4HJesV+ZWnhBRtUfzKue1Bvrm8AaHDBh5nMt+AftfegVM+fFIZEjOWaefcGXy
WNCKloZiSqFpBmPuQIn8sip3Ikcm6ydnyv1QClkyLj5lxC1CMZRrLOWMALrDyIdZ8OOeUip7+RC3
N3BeukqGU70+fk1IUG22jq8MP2JYYBUVzh3qamVn4iAiZ1SzGlK4u/vDLjC2/cBnMPHYSwIN8p4L
HPL84qPabCI7lUWU+1eSjvILE8ekYEW5S3VbfDSwQ/8LxAxtVu010fAiMmJ1ez5lqBzE3qy8M+DO
HtHbkGZdxhzFAziO+/R5uUGQBUGr9gzPIZw6JWxOMgLmnaaq7FOOPHGEXxf4/sCZl56TX+FvqBGb
RMBKPpGytcrIu04E/cc6ns4eWLfit4CqNUYYhZZR7FI0ln8oLLpbixkUgcTr3Ue5kZgk6ELUb3C7
ahwmEBOsM5kmAYI51dJxS82rfJN/6VVSMgOglQluoKv/QLGlIJ5yr7m20Fa+embA7JOglyAi3e/I
CYVtT1TJqJBnwueCipn7PHgZoTKMx5al3050lsK0uKcOc7V4/JSIhY1ufUfh5tM6fnssAGLW6f7T
Ul8/Dw9kWTwTSxDpa+x9cyHWRnGbvjurotRrHg55hy5C81HcG0QChczS9bGFbmv+RxqkW9YFnZ+2
Hc0mue2nd8jSlmUGFqRnc83ctxJ+lgcOFktvFx/gOE2GT63gcBS1YuzXbd1Qxima2wgWh5wgzuIv
KHuhpRRVgNk+STiLuOD/UCtIHay4++lpxPF4tM9yXyOkaeI5GkB7+FiK4u2DSyQLW9FkZeu6dt0I
AApcoD6I/oERqqcyuzqzQnCnwvSVSQoNCClNGnA7UOzLH3T4hOF7xm4GRdtM0boMq01qvyPmK5Wf
zOfS4f69//chng5ZGPCxGI90sABsVPb0AsQ8KhjvGovHjor/hSGUqaRgBQQ4ggYRyJ/iYZdJlg1+
pWa/aP1CMit7+pJ/33gQZYU+RxZkvLs4ft6eGwb55Q+GHvUr0Ix+p1nm5gAESzjRo3KF2NLPOom9
7DCfLnurhHGhuMTQ3ddDsRiyXNEqbM19vic4Ns02oq9ryQQBVyH2GHrVrX3k/s7ypbJjNzWVp/6W
o3aSOPPXl4JKGZymDTyood74zyZNTxr8E7kHvYGDSXTTaqVA+j7bzwBN98LxEiwc3bQxTSCJDuKc
yRQ6iJmdM4XVnGCPHPXM8g8VLW6vVyeqg5dQ6eMhsi7miTgtU7srpwz3DNSbaCcMeRWV7gPfmJ1A
+4Ot477fzDZpoeOZSR+hEe8QyH5GclyG7uQSpB96UXouDJOAa38rou0sOfu7/3Y/aHmB7hoF5zfm
cq5Lt9riiVKwp0FnjpWzsN9NBCAaKEa8i8QBqeM+sNRLvlNk9aqsntPhZiePGirPmqATrgx5oV0u
38KvDRaGDhgclx0nrsmheEY0BkpYJmIH89uJxs8Orax691D39Ic8yWpY9tfYOleMNnyf9VA1QsO9
HhOxoJyhLzS60dRb9HkdelEjDWTJkWpLsK0N6lPoevy0VRVGTbZRVjO7xN5mRIowkaZ3HW0oTH3F
zKCqZ9w9PRRqQitPpYsneCgEaxn0HjpiPo97Pxs2vEthQnqRiw8JRItPu0KMlBuFqK7gKFOrCGzA
LDYCZwymHmEAff4y25zQKnlQAh+Ht1b3H5VlWmlS4xiy7nrqEIPqJhl0pU4jztd7hzy53CE2QRNL
vUi8ovjI8HUTjMwjkE1I1OW2KgoSJZV5Ya8zIoQWBblkuQ7q67ASz39zn8FHYEbjMT503k+LOAox
38mRuUAnD0IUz7JvNNs1xsuifK3tiKcQkz+N0/owDfY6+vAjnJW1wqrP2blMp55/6sbKl638rZGj
o/aXFiWVDqpMNrXYnvGNxKfyMCCX9wk/if5ZpKqtC/RCMQTATX0V6OfUKAQZHFaWWFhKBtjo354C
jPeP+Dvlkf62+JOB7lvJKzd1Mp6Apk8Dqutg9O0YfF/e3mpMHrFl1FQazkYFXEJWlPYwNpv1jIkF
M94LhyWWIJ2kplEl45Mv7qPFSSr474sFiG1NA2Qw0NHy9fus/e0O1YGluAxFqalFS27lo4fTU+7u
kw5WoWh+ojJwPjXrrSsLGcAgGyywA0lNF3DGHuT3cJjWNkZInYgTAesUTz2jWZLof2IEmWm2C1hB
Zk/2vAYa3pI4tTKwNXFy6fr8vF5OYbIl6RDD86dh5JxH4bbSLtqd9mmOU9RNAaVSkjoM6XW63Jnt
R1ObXKVBq/L4FWILCbtIeepYsRYnIoxix1zzwQWO/RlksIaHjpwsZeBQdIip+o/1H6xyUTKg+EeW
8HBR5350d+8xuQNsLIt1B0j+jbk0Y5I/zB9LwqcurDfHHLup9kTmuHhv3u2CH8uopIUJk+WamTXw
2Yi0Ltae0loIcQIPqxcraJjbLal1P4ApTqGLpGp50sekYV0j1LWlyrUuLboSZ7rNj+Ql+U39jjL1
1IzuPF8wXnsioSo6jRfOmB3z2fcThM21xBvOPODdlVJIMBCFBMgstaJ5yMTubyde+ELDFkJki1TF
cwpIprNqOnvFr2Y/qrZDu4cLp9h6/fyQ67kozQEWWO7ZTUidWKP1gJdJgwZTKk/U37F4wSU9QA19
LOVQm8EDtH8VbcOiqnz6WnHOqvg7QbosWTmqSGn4LCjY01r1SfEYa8+0GBO8uNBPW3bB/U3klj68
e+yzxpU/0oKIhJUI4xfIpio7zc+kBzFSqZ11rvrCsAO3WzPMm+fjbsxEu8uxctpvYPycc1TLjBlc
HRhz3zGY5CMfJMpuLn1TyKicHJc8D+gOOW0zd5KvOpRmoBCXyjwTK2ckQGZORiChsLi5iq8i3xeh
GTDDkLOSP0nyuL2U+EbFHOu5mqxF09ffp7mZDtsA03TMToHyKC8WuqOqsXAbdFUARnuKw54dhNcH
7u5pxhfZW5P40Tx/HlbnBMcE1x0nGs1m4KQTtxjU++HAGvyZCCel8asoUDCgfo7/DvyiNlONho3I
DhPYAws4wtuPZ4UgSRyEbBDy7+dcx7IsAOMOCKkKdIo3l3JBn/NHGjwZy3dlat8WruVET0FnBJ9L
UUWF8khP6X5eneXNQi/ttxw5I9Xgsv6AgGMFleAghfvRiQ87j8ns/9DKVRIlJnC1iuwM7uVw4jD8
LVEiWtDCGx+qorFP7H+Dc6tCc12A2+OlcPljwqk/WImg+cr2KzUbYsuSLN7gvcNcaIJC7RG2e4kf
wwCvwJRrr0f5QL0CjEuW+oYNyzXbK0EA76/1Z5KGOVryf6FkQq9sQTzAtYEwK+Ttm/g4g30fsNhT
4F1vQ2s9DWUG0rCPUl1itQflAp9C4R4Zr6kF+Xzng0FSCNQDgqg5MohqCkEBUE7AB/Dk+r064K2d
Tyoakt/KguYy7OKmnSViw6v45jzaefL0Spo6HcG4SMr7ruKPbkSmTbRprbZfk49sYUOZptu0tXQ6
ASMypcCGlzZaJOKg20ljIV74ipkQV6Lv5v7VvWgXqAaemMVoUkD7JwV72lVdu7IukLdfoxYnWhrk
obOfvmp1jqikAS2JuRF2iRkdy7bT7IB35FS1yMktFgp6JlAhi6VKKPhgr82p5fLrp9pKsuffjq4v
AZTOOQAtNl/RbHn0rBdHJaZRz2VrnsFu0uXonOf8EGtLtVCPuOJuk/SiojqL/pCvOAFDuatDOMqQ
C5a63VCK5BOLhO0Gn8IIvBYuAGcSukO9IEESeDeK+Q2qDaE7Rtj6KfwT8VSQA6v7w1PgGTehddst
uGxxvZdK4Y9Oa9ceSlIQTiRGSUUI+iCM3jWZvDISB7XvofNWT0ClCZCkdlH4eRcTTQcD90Nxfqq2
ZQFPFoLMQnmg8Xw5Uc9OANohxsyiiXyYvGOsqXOBYmcUe0u7eGlQE7ghSlNG1yynELCwYfCCqJtU
VwCqMTk/6Xaf0KmS35fegrq2J1RSGrhFxtb6T6DGv9qR5Y4BCZd/3VRLEP8EhCzhQ3Ui5Uwmtx3E
AbbP4OziqtXYVwl/eeGEZl9Xx/QmEINuqjMJvEXEDweD/MmGV+bxWZJFWwQ/R1sz5rkC2RnMN4Zt
AkR7hwNakhQZmyvOI8nO2F/t9H9kqVpOO9CsZAu58QRYM0xQs3UHgj/tth1e4lxxaAoXqBcas4B1
m5WLoHoEG2pXBd7Z1vj0ynIqNlZHL9853BoPOiOPdoR7cTP2iSq4gSxUjQl76ROnS0dHTFwH6291
zRT4SNeyXP1l+1DKDTd/rmYf9UKwtSqPBmLZ+xEpRGCUA0GJAhrvxiJr5+KjD8Qlh5ZmSkX1mGuv
7n1w8nVPLfmqyuWtj8DEUTVES0kS62EtWgsTUExKLkp2zeJKEbUqG7LFnTFxC6/BXjD3cQLSbFwb
K4obgzkZtjFuGE7MM2t3bbq4FBz8PlcYLUj2MM5vw07P91PRgnSpZW89fHYBbdSO/lcIp9Nua5gZ
H0Q2SeQuj8fXWI6bJHbo0kwmoEBbyhG8iiKtVE5AHWa4Rh4abpp4XCeqC6gd0J6b1PlINFpPxZiv
KNDdeLwngZgR74x3z/oWyJebKDUmjwCBRR2jFSbDpPdWzgYnLnuPAv+z08heDUKNeOhvryPSaYd0
Yyjoa/C1tx3AXOchGX23S9Ewl1FiIuoTMbpJt9SEjj2mFjQwaE4J3GQxFaJgt2njI4EmGFrTm55j
+riSeS0xLVS2aUqQX2pD3co4yN8PdbkRq5MCBUfPWsMlXDCPGXtWG2gsKpi4Zveg56KRXG7ScsNF
SlwOgvEHAT0YIzl/94DPm+W+h5a3dweO0J1eoU/txlL31we1v3gvtMW1okhB+Mv4O96BXdZYGsIW
youMU9Jd6fpIO+tmu7R8F2DchFUBuxyHSBnG1sXufhIuILChllfCaJktk0q/NeFal7HZ2gwtKwQT
SMvYWEBGtPgRLWSC6aMJme8C3HLnurwTE6PcYjxRVymB1kzSXdtEUcxuLKH38V168kbmYwxZARNG
SPZ/Zx0THYpPFoh+LzhpZ1jpJNBQ0y4QjOnoG/FqE//VxC4WU4E6meg4DXLIXDpnAK6y+QQdH855
SJ4YGUIDZEAM0A8RrpYCUj5njtv2Skwj6zPrRueCv8BV7PCEICX6Qj+Gqs74DCkZv2lUUATeugKV
1mKvY9ps+prhP9PojA+SAdAZcFA+g6ngBTX8gsNlGfpBiuDrY/B92CbNthBijVabnN8kxyMWtq6n
Z1CQGXuKskTa7ACaQQpuqBEEI+YkpvSooJ2rgI+P8k0aUsW8KE6Tj2YsjUN8Q6x0E4eSYDgywya+
NwK/KMmkcmGzN526ej5bfR5JVLCaVZYZ/CDFjeOzALxO3pyNqxymi/JMg962MM7IJR2k3pEVrHuo
0J5I4shhGvfjVj8y71iMZdkqezqizqfT6FON7Z2rwAx/ncC31cUpDf1IE7pdb7hFh13f1cWF7eq4
OiMdTqtbkPZNiGj6wf3VZZLGQhRK8hBkqfDQz8ZlOAItGaQZl6VgnWrbQwZrepp1Xv3t5rVryzYn
0USIFrKDH5RyrFgy9/NkPu3L7Kz/+mMqrz7xDv0ezuhHYTmmR6d66i2TGPw9U74IlGbe2WETpF7K
fu/8JauhIGbN5TvFBHV7sCV1UuWex5tBA6gA+Tt02x3AbgpCknr2MfD4xrgkc4vW09bJ7zHhbFde
Mfhc/OBcR4eeLqKaaYf4+o8uZT4o6VoU4YbN66MuxMh52teBaO6LVapHKiXOQCAbhg4pBp30bEF0
Ly1xhEqOhtURazGa5TjJkFQ2puDfA0lvPEBD4J7G4tIvo9uG+4PFsTKvwWieZk9kt5qqWnklxVal
FNYJ9ny7+UvmU9qGFBZGlzcwZiVXY4cIwEu8T6WGTWk2rH+VDt15n/e4wOuafQL04SZhfZvI6I7V
dOwnt51I2DJG3D4uV4N1jl9ycftcRirFJTOlt0b7EjqYRme2yVLi+wgdT+bPmRYPjQsQBS9LVpqk
Q4jZD+vPKskh++42VbPMiQVNfBMTtCaetE0ZfABcpH8vz4aTtKzSocy1FIC+GhNLUFJJou4wMqg0
EzPUoVWwyVYTU2AeN4AAsxfJDC6IaRizXjhuruvaXaGeK91eUbpbmiN6VYOEMWd778BRryVhkhLP
niW76UxaVAaGpMBw1VSLj0gX1upHhmLzjWFMj8ov3W0XnStHVBPYJW0bhXIWNN5HsYvWvJNPincK
p+SQP3OH1E/vV8GiO1+zTXTWSFLg82xNhqOnbPQhvGbGbDz3kXU4dg5cjqae5HDIgcUjHq+2iTOi
ucEX3H05Z8HrCHlJWyNLdD5siTAl9+m2PcOY/ggLDU3UlZe0LiTVHSYuFmqy+uTZOcwh2UTZgBka
7YcM2FeaByw7sRMKa40t6WjdybHXn1yeDl6pwmkWzSsYcrzMZg9yhJ2Bu7+0sHGuXswWYG8hJxMj
fxSU4y/4MZcy0l9yk4wyaUd4PpXCkx9eeDpnFGDTH9uEpcPxIYrxjrB/qnJ08y71FochwmeGAE8e
+99zfqLZDyaPoz8iOwkzks+rfRrjoGrYM6bP4cwPep1LMfK08MJTrPjEvgNYD/piFsUui8e9j8uj
MNOZ4ziVMH1bOBKZGKkUeBYzwQRg9tdaZHTVaYp+FNyP4sDBRtCV3xx1XL80oBv2oldTSUk0l9jy
KtaQ//0u0gX/ZfCspq9645lm8mERYo9/Ep+0tSY52LX7D+TAPwxWORgHgoseQ+Maub89QQU+M6L+
5AxfiF1VSh1mPd98+I3EmkeXXXKc1eesjU95r+yzbgARbtAFy6Fl3gnUvZKm8aZAt34DbobSrQtP
7xiLYtVnQ/tS1EG3s0kq9DCIvnQNBbA/n8jTTLCvNcs9IWgcvDcroE//+XdvN09E9q5HBZx6bDMB
fZlIBpaujK523AvrRI3pDgUgoWAsEnlE/Lv0os8xJdkXmK988FxBKZk+Hu4H0uHtCDOzYDp2KLWo
LVoDyt8HMmLg/DmEO++eCLicJdDGwS2iY2nyBLN7B+xZ1apyR/jqsCQKjK3M7dKCYVsVTELrU7nk
eXrKT7ALBG9cIyIN4BjEYaMuhvoq6PQDWz289HUaxxqZiLzKwqQo2kAdVPBTaTCLFfcClcO0eS6r
DfyhC/3V9I3tQzCQUwgaGEjWzePQkCBZQiBgtj+Oktg8Idp2OfyKkFT/nwBc5do/AsK2WzM6umfg
Yi2hNVa/0N5HhFLAz0A+qmzpJI+1tMcKl0E4TVVrFtbYB1SAf9ywSg+Oq6ky+7wRqWCxGEjhhhhv
U72dNw6wKsBEvQAx5lOlKIjjpIh3j8ZaahlQ/mKesUGTeJPRI+MIa5aoaiSwz+710u7yaNJPCp9y
KuErX11aaNclytugJITgiW96sS97FchFYHLXvCSP511G3P73EBxkK4ZgcgTsByKsb0lQ5ST9V6fb
vEWOwm/MTwgYpy5mFtbCURewGHFMF+oIMPQ5RK3LdS8uEPB0ssao66/KsWBo4SC07mIW5Zvni/3Y
xJQlItSyAt0ODAKzpfAPFyfbX3q/HDpu9yfY1TWjge4FFZQ9gA6+oZTiljm/6ynJv/xnU3Sq8MfJ
APH2837npEvRr5wsGG+4WH3Wh5zkxuuOcWH4JsDCdpKImfw83jjVx6ALnia2JZ9YcadYI66xHHfE
wLdtLlMjsAftOSii7GXZSfSiS5jj9xcdPpxZttPQjdFhUK65adDDH1yEsapjehn2L+k12hTLlrPu
H9w9w3gJDsE/leq9vvZCOUa0APldlXW3NjmKT4M8uShlxtuSAsSuwMptIBEg4tvu8BAX7bnSlk2Y
cWWzQJSPhDQTv3ajiuAvewqd5AmEQaLL/naiurptNi8FHmlauk1IzFcYnqThxRMljedKaJUt7H4i
yKV6kSGBejhOKW5S8S0s+UkPNWl3RTlMcX8dVgT/QoahPqx6mkG8ihGWIXU+1AUezB3+jRtkUbFr
ytfuc9rkrMJUMEjI1kfXYE40pd34tJcXCslZmWFY/oU47O7ZXpCnQuBoO/32P6s7ilmilLBHsh8/
YFWAfpTQgPYA8D1A3jmTVqigN6CvScsmpwKji1uAQD5Q8yCVO+Y14Ju3Q3KB8RLwqjdA5t/8FmQt
2tmzybpIgp5VyPQwNHlzAEQwhPDbwb4Y/sy6aPAs5S59qDQo6gY/55oSZbnIpdb+GuSP+CwMki86
15JpSkAC/FYjTaMwoAwUTaHfDf8jvlvAwEyXmPxKb9idK1fPJCXCOfwuSTAxG6h5b8ornmSYZFzp
DuBhqvHNut/eAqqEo5eMS3xwPtkcnMRlN2cutGjUiObMQ4oXH2KjHgq2GgVTH0ktlsTYTykxoyUX
F49DHN49zd40oYp/G05wc0Pv/Y5lqirG0gzlyUfh3kfPpbAy91hDxHyWbbNHHMEawx0I1llXriNq
21OOcgxZcQpjjAg9Mhfipe2z4M33IzvvHKtyBiRffyrZvNonOSXfvOq4VE0ygqcEZHLt0uoM3V5u
MkJAtf3EZeMgsuyHy4mavMg2/MAQlpR+QvSoeLXfEaQ1SscVE6fEmLVwLwg6WY3iYkfa5HYqHO8z
DUnnr8WyojqsSQT/+jbv5uVtKSzVxAPCc57eHU6pty92D1APdMtdOaHfql9Eb+yMaIq53aw3puxD
S830svfiPqc54bwwJBsiJWQG0ULNHKjcHZ7gECGVHxPWjwPSURAwLIGk35BKm4rUx9rPspU3I7y2
a7k077Q3hC8pqYHrGWA1jGeeli/+W0D5EI2lvOivks98SRSpNiw7qxtTp3DmeA9SVs00RFXUoTGx
Wy1JdfAesxfh4g7MU6gkI4UxVJZseLykfitoXxnoGSROc9IhQ82cLU24FfoQ1AkLj2SywCaelJ9u
XpUij5ai1TeQwaKVOo16UaCAvi/BBK21GVj8/AS7AYUk8wbNeToebfcKMHatUgRpXjZ6BQr9E39O
5cQq5hJGxN3dEiI9tBuNAMVcp27gAF+tVAUog8XHxnuePC8E7in7Erfpnvz24GAgf4ZO1ELTN4wv
M/7Eu49TMWFT5HuhGZLTvbpw3+3kGePiHgZTAFO7a7Y831en3orGLlZygJ3FXT/7emblSd7gnzxB
VIdMcUzsuDaZRr10HO8eqkhnKzM570q98e+Vs+1VEAFsSnbzHDqefKhRTs+anLv/QAJOXDcN+ZzY
1gCtkWoqwltAdPm9Ph9dT813dLT86fHRgltL+zhT0c0Ap38Unu8jDGPJyMzq6N8qixOXd0TzahHB
y9KS4dl/b56o0t7cjyTIvrPd3jqfWEyUnEfVFRqnnNQliK7CEov4ObvPzPoD51CLZWANQA+NZui7
WWzQeKLzhwck6Rl8tovGGW1TuQT/tdWuyKgtNlhjMTRihg3WtS5hvxUuB+OEziy4rhhPi4z1pEI/
AiN2rhRgu72bUa4hO87d1KHBLscWS/D93afL67+ih5cCwRDjUZAzO9a+TmWKG2eYJ5uBXwRxsl3L
iYHuiQHiGbJoFJ1/Q+vyVZX1IhRdSwG7aCGVWNcPTM2NuGj61UfMvNIFnWzEdG3ER8QD98s3i0L0
MXkSBg+CjdITrpxfU3cWBdezesEXT0fyEsw9DquFVZSRUAgt9Kzs+5PYgNpvB/dE0eNd8CT2pWnI
d1yQjQ3qLBVR27Pl8NClC3dM7upGuOjH7I4BRwnlGCn4pwLKdEDtkCBHHvFEydd0SfZiPFts8nYG
N8J03X3JmOX1eyI0S8sahhxokx55k/5P6HHNnJFHT4BmQNEwCL3kvajmGf0eCwq3B53h/5zTQ1Of
QC/S2TL44wW4FkUM0qzc0wGLyzPDmsXKuPf1jXA3ZVeeXPssEp/5xF1T2S0JW+mU4LSDQ0dGGWiM
/rlSocc2WunQnqFbuer3G2plYxGWdwMyFwXfSRwJm7pW/iPmdVvVHZnisR+K0QABWmMszAPuTvC2
zCN2KMlOcgXs6mSX806Mz2QYcQEdTxgJ3YjZGcmuwicrXGPYbRserewebLYZvs9pgxmVvTYDuKYF
/GOqWTblAKYFId1w1FF7+HfJrCc1NLvhy9nSBAGK+k4FPaH2Cr13/tr0XyDDWxMu47QaPxHgTJ9d
uQ0ckeAGavhpA+bZT03GFbzIFuzn0eR0v2Kql3+UmCNhiHzD0eQiAnVBLg71NM07J5DfpagxBRqW
Q7zrIWXvKbCFALlgk9014b7j83v3DJ5VeUM2lkc+iV732R65un0YJ/JWJAhzc3h0dJu6o3dvxHmq
GE0TSG/zdFOVaFUvQRsdcDG1z+I43n/XHv7arFnV9mVOZvqDPPJh3vQkq191jvw3V6rEGOAPhezq
k68KmTjxwpDJXOt14Whfp0aUV6HMcbhSAW4o2b/vGqSqjkLht65pqcgCnjZarpYY0+/MnpFr5XvO
plsSrmxyT2Fwrf0D7b7Mqj+/fOjj9gOFSFSmDJSPDlubDr3jT4yjvg8jIA+F+kZjjEaVTfjSesNy
B3eYxYw5hSxOLnNSpEGAeA2jlzv1jRSwmH+roZArtViy1Hwr5n/l5veN2yrLEELAsBfNBxtl46VA
KjHsGP6ciTUi+hhULzoRwMbY01Yz3ycmfq08BT/MYoxGjr+nRLy/ZL48llOsHveRjjP9UHLkoiL2
xZNT5KuRMpmtGmERijCTo47faGIstdNMSNAtORd9LlQfVMzfWQctHXEdyHkC/u0S6Qa3amaHn41m
q8FBsDBl78/dUVjxEHdxBtwv54Ys8AxDjTsP77FvmKkVyoKWL3hGBMgfeX/US3/0hhXhVJo9+9f3
8Qy1jwKwn9UCX/Lh1kllVdSOL7qdKfXIW9sW8vWV8dxkZ4YICtEBzJIbc5ba/xjso5nFaKC6j6Pi
0CzQBS4UEdE5RCMtZGp8gCY5jq6uEHzmtJcEd7PBzMXn6Lt9V+MIJHn9WY16Dkm8HvQPsT73RlCs
TfFuoPi372p/m8gCrXUhwfLm2GNTAL6yWaJa8hZwoEwr9vkhcHPpaOP3atTz88H+4T8Kw/Z16QWd
ZhsPwvcjF5bVlrE+aHh5NxnG6S5mVYW9YLYItPhDvY/E24352whwKSf4ftThFHi7GDNyq3w9Dnz8
H5l4O8YJLhDyrhTT2EvmqgWMroTTGXNlMV433zpAXBBnWJ9UNPr5Y1pFW+ZeDLzmbh2EtMspNNOw
rSP4e2o3QnTTmxQr4u3J3RyFDMrbpob3dRN23f8y0bbbuQuHgJd+5nBp5OEAFZ78aRD9DAHAFY+W
y6gsqEOjvUQ+jLwDXoY4XbStR27bCPTuh0R1WXNjc8OerYwsDTxwGWxCxnvXxae5c0bP1x8HHB1A
mG2JL++1/Ja8pgcSk38sGKEObwZoOwqlBC7E3mR/CerxLLBeuQmfmDw8hKQ5I/rgAAgW7JrWK2gc
8jjajfjzRh3YNIaEHJlEGtzws1Ch8GQiErIjQmAveICekHYsYhV4a4FVkkuJk5oJnBvOH4y/NmzW
RfBcntmqYkKYcPXJnhFdLpIqBjV34YXEXjd8K9uIJkaH0LEJKBn6soFcFmujBPlpH181E+XBHWyE
EEiCf/QGEs6dzXwPzPmwC3AeZaCY86VWM1y/HfIHBn3yJj88+GdUsCmv7Tv4vQYwOD/E2EayYrc2
cbqjP7CPw6Bd/5mtPbOmaj/MNxPFrEWtgsWwv/C3KVIjBeW6mGxeU9rGLQ+vrweMuifg8hsPz8s5
z6G5FjtP9Ftk2exOfVw4ZUi3rZQclsiHE4kxwRbWHLdWBM9VsR5aw4QGfA6LBxjHvj8EQe13+fcr
7Q/Wv83x5Y/+GYAIKJKDsOWbvcmTs3GoiyL0jGLNEMus70nV59gpK6DwRRPj7lztgkZ70dxjVi+R
G2CucEIyFU4jQWjL3if9NruyuKOiUfVoboWVjSlA7RaHtyvV6ZAYpd1JN8XEfjxrRlzL9asuS4gW
y2vxtW74sobuU65OzBp7Xqpeqy8huSDzqAtYJv38S7doHsnENxxhrvNcqCW0CZhF2zX/0sYV419H
5EQUH2i2ZJt/riYqxWv6Xn77icJYTLHYGSososCLab+wd6aPIOhNxv7gE/IAtRPLEpXXVk/ZFPkN
442JvAIeqfyaMOEBa9LHbNggiVw2BMOxA0ZpzECuLiuILqvhw2wHRrACdKHFc563EdPA50xyNpT4
QB20wF+m/p4s41KZCdxGqdGJikeJG8RbUiYLnXTaDsBLzA4HiLVjSSk9KAIlvLWzllYtRCXBKrOt
NJwUSSfXWPeKisKYLjfqV0D6pLLhqfDS7Yodo/kObIIKXLL9JFXdt+zg0W/h6SgPt4GQfZEVFzEA
Sn7A+CSSluss0KHmrw7Zd11c2Nku7/qZ5sSl6o39H4GGyLRCy5CxLcxVPWoGt6Hh0vZuChdqkErB
duul6xR278LmdB/3kD7jPrzVz+g8tDlUe5FWezg48UozkGK0OA27DP7Rw8+k43NNdxdz6MzXv9E8
d4ItZLTlqFIIHrYmxQe/1ztQ0henUn0aLf67HnOt0Om5gbr909DAOE1YXfj8qnsNoU/UcuuKyTrB
213/Q1eFJdndGiMuhOqDP6SR9xptXMBMdkwkCxfRue5LBleyo/s9SrlyjDlizJBI/te5MriLpwZf
y6Ok60r/4U7R8BTUPuf/f/8oNWlG0C5AWfA+EiNPxV7g03m4Mkk41EwDJnwnmfwKAMpMYszVFhMv
iwMYDH8fpOM+SRie59MConuxw4V3jTBSMqmkv4g/FkxUr3XHxeKKS0Zefn1XtiK369B/LB5gM26F
uzqHiNmjY8xT1ugJsyjujemRhoa4ABAS/WIivxmkpZ2ru/Z/SoHgf5FhHvn0Dk64UGzwhpcEOKO6
5HZ63lnpElUXN7y6WIzbECMB2U6KCkOJ7H+kzLqJH+sVQbGIAjOzQ9eyHniCARsJS63cwqIDl3ld
R0T3P4t5cq7DTIx1/WcLqXW9mmxsFJLUEItn9wQE/kA+TA5KxhcY9xgTzqi1ifFtZQDtPW428my4
nRbriDfqWbLCqRmzvHk/OsbwWeO53gHIKYn1xpZWB1g1zdsD5ACBpEgagjfSJMqXnUysRl8uy4mp
o8XKutTE9BRlZQtLHrSZkU0tJndduYrkmvQM9zIjAhNfNhYql0+6P00YsaOMyx4ednkC6Iy2qYfN
Tta1NatTdcxJV6Depmo3ebRzfjZDgb88fFUqXB593ch8Xf7FH5X5MHb9S6eQuOiRP+lFFPpuwZL2
Vl7deMCokWOU6pt8jnWgEXOZl8jWXUyxfqO12gu7SfZrDX8fvEn5boh1HrXXJmvZG0rT8bEJHnYi
MJFX4T1zFOA/IiEFlprGbMUTItFGsM3ApDQtRsIn5GqNWBOXYnc39sDGyr7d4SHFEFhfqBcJMSFN
YbM6N47iQNPUYhS8LqU0MTuRbL+gpyfyotMLePSR6oSkn5c7Sope4sEyEiuJWbAXEEtL03FNqjyo
9jubqPPyMH7zEOifX77IvclB8kDc1XsAUjhFVZKBZace4lrrEA4vlvfYyOkZJBfKyYI71oiC5oIO
cYkbZ+b4jJaX0r3rc/wxHV/+pQGCTXbli615eAGQhKYXHjVpjGJVfCHnF7uDzUgMELPrTheu7EPM
tobzv7Owxquf68SWPJ9eHRhZ9nitk2baz8zMD1gNML4kGDwXeHSjUs2Q9XT1W5lkQ3VF5J8C/X6I
syxkDLkwsADmDejlW8LvY7yKnaO8hYNvWUEBQzvJ5n0a/qCduai+VY/wECiVLwv/G3sz6LaHea9K
lR58/T8ZJnS+ouWWjWNfBIWLiNMVyV8XGi0QZTSHVwe9811Vil/722c4NLnzJ/wLn/KMtcwdGN5r
/yCwoLA1L9wiaxgxUyUuXg/8IWF1rsxlQolucRa3vv8ZVgJtv4BDDqqSgnax0FUvAzeZM+ggg4KQ
nl1ZwS7tyO679ekGUCs57P+WiRZSDaUEhdHsxLZgv2TR5Oxul2Ig55ml1Rp9+iGPh/IoM8I5ZcLp
3g91re6eKPNtjNyuaEtnwOq96/ym/m+NxCz7u+LE8UTqWChY0kNZ+kP4LXXfaus8ES2hoOEs+THr
04hAm+bJbrvQrD/2PatgGrUF/0aI8cdo3gLczjh/tNulaDvaXJbFWG7FZkOm+eDfQeTOvNFgiE3G
54YoIPq1yKixlIF/8bAHsPiVJiGN4MeF8qmvd9i5wxVQwGhWziWFmJgjbECEkffhISBxHsuqyl3n
bDVoAAv4dzR3cQ8MLDCZb17KF13GVqJ1cUW9dRlQuhQRlfS0/+pXxz4sApw+scgWHmj9tXXqB1GX
DHdaNK52nDZ7pWuq2ol5htX8VMz7iZkchPTX2Pr6y3lgT1lBrhVL08uOsWizPjdSSBa7SX/4+plG
/8tx0VS27vMCn49YZEpsi8nqz+Gyx3PXqKV6wHASCqlNvE0f4PTocWpk20xrqxHS4PoMCThFSpVA
xbFEhG2EZJByjI6vD25ikKNCk2+YiTVwiG/mDRKMS/Wm92W8MEjuQmOdSiTbPGe995D/RI3reRP+
BN56c6EXmXhNlsbm9Okj+CdqMC30kB+SgroCQHSfsRrUVdTl+ifU70qbuEGM6lFerVlaGHFkW/ms
SlulOxFA+Zgzphr69JWdIWk6Pa41MdaH22leNkuX374jcjPFvTFt6MXVoBb1r7Ubv3vLDmOp2lrP
f2SpdWx/Mfirpu69jorawrYyG8WziO2TplUPaqFmASpzb9DXCgfg0DLlzshO5r7krO/6sgHVj8rO
Bzsgr5+eCJgNWkVYvG51fg3VFEBU4tH2QYA6KFKUyeQ7a0i0CnLNU6YiV98VAkVFzEF3W/J1fyld
w+AjUoTl2U/e2wnu4lv2CxsGzXTUw9gVF5Rem+UbVocHQlpzrEvkh/iHXhJZZOtpJQILMyAIvQMt
Kc4adHYww+bNpIU0Zi5CZ+NkLgB/g9Vmj+TKZduXvA4S1SWyk1TzHKPFWwaXeq1zLZ12oH5VzjMx
pPUn/9vS7CaGihSW2ldaTOAqA9EoVVE2AF3vZXVchRUHEYR992muDrS7Knk7J5uLZ2Ic+6iFludh
9gOzk6lLqopD44Ph5DUby+K4V+GfVIgW9LBvS+7HtGjE3aYYbANp9wxyWUzPdTIUNgM+D+Eo1iXy
sFvDESlVhrYTzUDHpa/IbUUAwptV6vK+RooZyg0zLwGItih/pvJ3P3UFS3BjpUbNtZJUVwCLhtWQ
vzPd9SpgEyHZexiz0A0sfjrFYSqeEJUrAraHj8XlfdSor1eFJ6uG1GHvoLgm8mbfbR6W2CfQLvaz
+l7Bp+BzK6rMIFFS42xQkJVz3HvtwoxeLTun5k2WNvg63vXMOFwLp8RGGUwbntgi7s9MlEmcLuHZ
GBbpd9/Mn6xT2x3YHMHVP5dzt6FyMyf3xda6y1Dl12xcaj0kxPqB4GlPaHgJfm+Ie54Oe3wzYChW
0zsxWJc/CxSfD/lxUxY2Fr+70Ze04e8wLJgaiAjlMA2j1zII3bUf4Da1YGxCFG6JmQ/Cqx+LRv5D
yKrk5uklStMROJxFcl32biyJ5Q1IUgg6PHGo7GJIc10kQGk9QboUefDwo/TIdynrciQp1+TlVzua
Jud6Jq8q9VlfQAqrmoMogFKkh3Y41wnDxoIhKne0wofVoOq9MlGpZ91r+YKUIOFI9LfOLEnC2fdu
GKbePXZgX8VGr+wUmYxlmGj+MD4F+Kb592NoCBslMuxRAxjtAoN1epIlohDSqa9q1M4V2DvXyYTM
4Dlahzgb8/f+30DqH9sRWAzcBhrDGCE0EGcIulZtazvS/dEt31FP0mZDJ6POy+M2G+AF4cxK3gln
VeruiI5lMGoXBISBUMBXhWtjDpgV3IKZoC0gYPFv0/lKN7XCMBhl4RzBOudoT8BtTGsxM7y/r79E
mZbPH0BE4MH9ap8BWUfgvP2UZrVv3x5KEoScabDmh3DLQyEscAEaiEKmV3xGvWedQkF8mGUhEIAL
ihROH4bRng04o7JHq0uuzjuH+uwxh2XaJG76osF8KFNbM7gBw91RDRf0nmsU/jIZfUUO7thILg5d
TzB5LMMvoZP5Y/iakML95IfI5yktIPEaNaEFt/i6KHb9235d9gauxJZ4mkGvqZuukkelbi40Zswf
dgGIh4JWRWsV2nOddGFaiqks6lEXMnuuWAaZ8hjANh+ZJst/UdCDER0hX3iR4FK7gxqRW0Crf+ja
RfmOdF3mEkR2PZsJwMSt0GiWeh7wI+ou9DuJcEcfheN2dMpAW08VfOgaoXEpmA1i1UufalT2Chgi
z6jyrVWxby3wyz5X6c0QG+9ug9QRCEXDEdFAkyysZJKvWO4U8JG1ngY6OornJv3VFjpOOnjtg6pn
ZHCi9wlr/WwyCqLIdIsMUSf8MwR2IUwXaaUfBfFbw0akigVOA+Xy6zE05UCE7yPb9TIfDuHu2Oiv
H+h2br+E0w7sJ7Xdr7ei5BgwIRm055U1V00kq8naEOSYKrU9J/yo2mN359HEiqRjHlCVkqiEi0WD
5DfX3Zd6HfAeyGOXI6akLMuoIkgRSbB+qNjsbUTW9WYq2cYXUYnWKJ1IWT95csPPMU/XOXSv4Nzn
39pc/LnSAN3p4jMJ8aVCKRNFFIJs9QG/oRDrz+8kmIm/9QFH+m9rhoRKQtV/s2xEl169XYbckDJ5
1Swn6F3vqAD2u5LTfo6ZBqhXHwZNqrr+Opnsf9tBgBJtDlK1h0WFxJnFT5e9uMYNTv8Fg9tjuO16
HezwLvX18wN5zrhZsPNywkVXjd1ZWeR2YlNJGTI3JK9i11pej4lKgJxNGKXdFut7hF0OrJEFyPQm
uj/tQLxb+3pt7ACHai7UAPGzSIYnSBl70qcrHGAxaRZApsGfajkpLep6oUfK9jnE8LrZVgEAzD+V
KvDOxqrol36P4sDQnZvof6FtsMEki2MRtLoqeE/q4GaD7YOX0cZ0vCyIoxvSIH2CFQUvvAGsDBGn
2DnK8PjCYQSR/5B2RKL0yfPHJ48cO4r27Ybjv0WfbR8L/D/rQUmknMMnkUccJyLL4uVUWyEdpw+Q
2k0Yo4KkFXVg0nhDC1xH9yqhPhzn+FnRa+c4M3sxvzCaeM3ja8aAbmXBjZjo8u9T6DsD8JF4hvf+
+CNSS7TfngMuzfx5tdWhRkBGaGG69JyAtKBeZSggDWT9ipmh/9G8EsVukcs2l2MzAU+X0IL6rUhU
G8509qJzD0RSXK3C+CfPF/JSc1Hwqkiaq6ASgaZ8srnLEXWX+gvfjHPCSuw2cJmxWMkuzpuwrZ12
uAzVlSqoiL+Qn5NfShO9SyXytqTCADrg/fHk0UFKbXVqJT1TdkaYIsMPs2bcN9YfXkDcS/42TQaD
URRZNmuOIW3Q47Ed7xmzZesMUq+v5opMnGoWUO3ilak1/udqQEW610kyjZmgLWfnNNMjVKgW2jot
djcLsRr3eTVjlgK/gY050kXqVqUg3pItqRjN94LyDQXccrNZCZz/ulUVkm1WFBztjeN7vr8tep37
Su6BdGxjYVJguduyTxxrL+tYUoiiP7Z3WGlRcZxabSZeYJtbeFDCO8LY8KIuWUPh2JSCDjHzJONk
PnEtxBXDs78HhVPSUSw+yBpIruJPeP58jP1bjPlRoKed9CkKwSZSNs3nOo1PrQdmUhXqYv1dTnR7
/uh3SAlIUT/aKp/BVBGJzUyBm2McdSp3dnOoJtKrqMbOX7JzYUuqVhlvt+6Uw4IFdwMO07LiKt8o
OARcjWfsa5UCJU6ojRXSJqbgNKAl3JSez5k0+aeijtjbjatv6hpcrqBt3Z9/cvNSJ+ZNZysNNYDM
Prl5xh5gIYFGo7U1xyZIP9sVCdzWbtVmGsTCu+D1MJMGwx6wJKwKfQ8SppjMgr9m4rhrE2RV+37z
6GU5aVWit8yAV394CRwgMRjkBBLxVEQqteEU0ImvS6siUpG2UEPKMXSb2xXnDnecsVf/g2iD9BVi
x/KlPUxHpC1eTr+/O70EtdbT+0c37X7rlZ47AmbcnSobRhh3U2UTn7qGtELbayvYwc6abwSoB+av
2Jm3dGOdetZW5hhOObgkmAiQRh+C8d7XUjRTyx7AT92bJ8q/RiL/kgCvn69c4puq1Xvl0a/RvYJZ
JR5VjggF5RzVZzqTigq384bjHvwsxpcSWfc6TCIuF4Qu5mEjx/C+DQAYIbfzVkvTmZlBcyMxzjyF
NSx7U2+QaZJA50w7lDdbdQ9WWbU46SnipJabS1JOO60c/ry9GY6Q6qRDp9evpDqjDHAQO8VL+SrY
LcZVpwPx3Sz9TXz3FRk4piu5fAkDRJlDm1mYBsgNo5p99eGtLn1KauB5T2OIPZaqLqLBYk+52TmB
OuBFR5fgN6gOrKk4tj2FwpJ03z5/UYxGvp9XBZGZXmTwE40GtMAb2HJ/NZoODS9cacFhhyVlOT6f
yL2YSKg5nBSWqwrd1s/XfcMbexjYvY/kiu41ZNrCM5wlMOAlAf4WLR/gb3kjEf3Nb9/oMwoszXWj
w5chkt+xpu7hj0u3Ia2k0msVAEAkaUyPUr5qZLTF19BecMIL6YfHR+sLKihYRNO1/RAnajUq2K3R
hXCb8hkdx3qIJ+Ymeo8Vbxmb0lI9kSdR5IuAIr0nJq2s6EIs8MB3s6ZghjTlt5FoPwDI/h2a+Bpg
s0qEvLpsU2mR7T3PiFSWqehzYJYN55426Q2cocamqqEls/ygL71Vqfio8hw8Vi7RkqiyEc45ImK+
li3B7R2W843eGWoqrAhpDYOyLseXzHpFR/xO9D21ia9yqFhq+GNCwzEsJT3TvX8R4X9Rkv0zQ0Sh
zZi7krVN/ro3LQFKZMc9k3AH1/EzFPnhmNV6ZMvlZknk6ItKDWpwNxdaIvghPGNEXl7rQJXX0Hau
T+CUBSNZU9ajU+wT8C4WVqyp+WRAaUjfpDXo4ktdUnn0DOSCPMvs6eB0FnduHuShOuxXzDVp82rC
occTU5FbMTXCAMIKVPCzsAk/nXdxSIXK+6N9yjWIduPb1AW29ec60ZrXF2e0gpglR4nH3yzd+PEQ
nSnwnvl0Ct1qbrxDLPv6HLDnEPYkR/Ln9csAmoa8ks7cl0oEIRnXjDfKng3urW92jVsqG3Sr0vGS
QdOe0gBwEsuPW11uAVIQimnNYbL5UNC2pohMQY640HUTSRV2wDdlpPF4a582H9SW/g9nFmAZl1s2
UoeNPHNpnMz5c78qR2mwUOh0nRHtZ6+a4qRWQQLk4wtBfRBWQwDRTOjIipGc25bEQ4KIH+pbwAgJ
pEkjePN2af+MfUIgPGxCRNZrP7aAv/2s5+otSAGGsChakafHZthiBa2SZcVfZbPY24PTmML6gayP
uhFdur2AOuCQY+WRLDMyZhqe38KjUkYpifHL3w2ieiWPYVDKPNXAlA80QFQVxNFs3FfKyU3DMFEm
6abXv6b/fuTAbWQgy/wfe7Z8/CAs8PhP6PBZ7EmHRnsN8ODN6YKLb0LA6/5XaCQmBjoRwOnRC6Xk
RV0V5qqBaWNNCRM4rWT4nHM4Rf4ImwgBZ/8HCiGHiCDlEUZi6Kbot8EaGDqW+fKlFcbbZGeBtt31
S3yi42W4d/XDNTJjZpmGiOPVpDwjtOoMzeD10twru1Pqj0dJfx8VuvCEMrLL7rJnLt9wHfM++MlC
xFBd7UNhIverDFn6lrDza/jVcvyxtQCqpEldNbXKAsbXo7CcUukJx4nuX1PtVEACabCXarVnXHxg
sx8T+tyVr8ma6h6cB2OdcnAQ8T+a7kjXDR17lmX4p2sC7nXdWnfB0fGVE3ATbxDLdUP0h9jkyjF6
OmoR+e3EKVKmn6HXXWpblVQB7MsOrETokG/C8q640FaK885VQtaJqktkmcg5dsceWCl+5zST+/uq
S3vXcuMTJadZSl92ocMhtXISEU9dCN7wq39Zx+EIGWyvPRSupwEK7Fe/5jLxPYSGymcYr4lkOtgx
SkR3O+QgW3ejUeZo05DbmIC6UKuE7Pu/pagZc0O5wIOwqLPuCbkTrKj8diD+MIvz+wn/10e2X1jF
L7duHvlDyg2ov9Webn+EfE50qNHLgBjCYGTHqyQTNDfI7iAadpUFrtKdYljaIBjEeQ5sASC+T53l
5KwWtGk3Twld0E5iB2gLlTCxBRK3+Q9MwYxEuNeAMtT06uWLGubchw3otQnEiXX0jYl6TniRAeJA
MeVlG+EasYNbdAxWjpXkRjQXwPlNfkHCt79YvRAvE55SKRACI8Qky24nea7Xp03oNL4jbwKbW3HJ
KRdjs1H0CFnBulT+2uEnTl8hHH5uHwG0ht3oh8KKaWjBX7gGZjLT6lIDTRIb3D6RyIP8z7EdY9al
SdgnLhK8t2WLLIVODyspuv+vfGxvVmlgR4xwZqVoWHrYhFoubm4qFwjdBefykOtNMR90N8QjmTrM
oHIsQ1qN8r8z+Hijnl8+t6k4s15H8BpNPVde7E5tWaHVCGc6JV0WeJT9eZzhw8YQepsw0cmfhI9F
HnMuQjVIsbpqf81yVpP4ZeV/aaJ4VYm92zWW4J1/Ofh1eL+ojd60JwOJuF8WmqhqhwjXjs48FZVn
9NOepQueQQUWlccJfiqyYOitumrJZisJXpNwC6yGOZQi5ygQQY4HV9TgsbmShCSKxXe5GrA36cL+
DMCZ3J69k5VJZ2H8WDVDvZ9J1pDDh+ctQWst5TVYq6ZhEAyAHNlSITtI0iUH2OMTCIyNAtdcSh2m
l/0JwCyp++i3d3SQl0xEjkJ4Ti6PGs8wek0MEUdiSaREbc66LeZTm7qZnV32I4IHAg7wQjCCKjjO
+/3h0f+2GkhtbYOvyl5quh6bphdHj5ylZd+q6X/4sEiQURU1FscmVReFOZwtaWjHHPVkZpTAFI+O
5Z2cY+WN/wL86BH05caBncCScVHATQzEx2+txaHeGXp4k8IlM1k/tWWTFUyRWgdVGzSgCFASXLz/
T14vNvj2/OowYOuIkdf0hd0Z6fJ8lXqU+fMNQdA8WfoQEWBzurwOQKw+s/nR4lwbbKIXV0l9n1OC
LJ7RhkJySWZ1oLr/lVENBO6Tdb27ErARMaQ/OfoEp96LjrisqEqFe/ByWxdml71eFcGcFsKLaS9g
astDRMl3mQAgCBrptLhJDlt1khITT50U2lqhBqjurG3oXRKLyTOXVBeuPEdlPmyDzWiN4XOtN8k3
A7S2d5eAB7Ud368NDnyviElHvpyGJElWYNQVKBtWL16DvjfFkqE8INYzvpf5lc2TWsbRHSOnSxZW
O85+whO5MmmgMCIg1YbTXc1ZYDygm9Od4jIMtGCISKS0yNEa2uPql3aZpzz83IXvSherj9weMS+4
TNCy8VfDudBwCZWkBNX69wrzVdtWutsTQ7dhG138KXDak+tEiONFuYa4FXRyP44E5ZjTZy2OIuFK
uJPK2LLKDYUsTHDQUyCGfE19t0Chh2U34ExpJdSM11Y5VnWsRxtY1epGpXNVpupUJHp0UUgyqFJ7
2jhqEiGQ4Xj8vDDGm5ePSgkiwbvp681lBywC/wCA3Ux0nA7B6aH11yWV4eg/y90hj17W8Cx5ZyJO
tDd5KUHU/085GRYDOHkJ/Uc14iFIRv0xLAef2Fs5aXrre0XyUbmHhAblykVvjF74oypFLoBkhWIW
EWgHhU2UHRFe/DyXpAjyYuNJIKRA2eCqVvcGaqJD7yuMIq7TMBcK8i/URUjbjkjkDmfaoU5hcEM3
xYdx7nBzqY/Zq/v3Decizx8k7OCM33KeKqOMEhrKUaDmYfxMAmytiqnp6ycPmVtJMzhaKIs3KZV0
uKLfYz3sUSqHsyw00YfqaXp4yl28auKmsvD9skHnmBm8XiyBweQDwxaT3ZCSkN/L9sJYNpMX6jUN
fcyIVfuwVNByl2TUbwzDinS7+Nz4lxGv2sb/eP1xwN6tDq1E3z5Ee9MSac+OTTVzOW3mxM7LCcW3
TBWzqquhHT9xYMjP53GXTkLFLJmuMSCCSdCTrjXPtCTGc5SYUHqVh8SsS7SHWFMv27RepwxDHYys
eSp49P+p0AjjtfX3C9CSsxjgVWDw94VWJ9hvsFMuES1jWO0MZl5mvPVerwLBY/qGXiQwVfQjpOCw
46lHtqdetwHHjFYUSU0qih3aLQRdvsHM95olMYtG1FOhHi65nb1/WVe2XVl/aVCOLrEOJ0LjVIcY
ZXbL6Q40z4yDzOIyONrulwcqUdyAponpCKyaY8MlOCwz/ESJOwhOAI/wXBLGJ3i0uEphKk9mS23o
UjethuQrpi/OD5jm+gzTVs+UBI/rc+GExyQeMlqwcqxA8HeQgyTzaDF667fFVrEFDackfxe6ctj8
1VFSfbHrJnOHCfdbjhoOpJ8Dy4ZXy3FbI/Lkiil796XiRXs5r00wdZFsgzTNtzF6VURxdsDnKs3H
9BjVAvavV/uiD+pylaqBzPn8WdW96IWC29x9BX9uhFdizlr3BuSQmamIXE4fYk9GJYU/+JUIASBx
sbKzQccn8QXCoASwWdnvDdBvrEjJD16aACITVwQyG+eqwRPF9dSxe+onGli/zcD3heUaGs17bBes
QaSAGF5fXfDsU5Su7Q7NUxFIUs0CnZgKGWrq8bD9elCDYmd7qAtWd6n89Veo60owK86DsZ+r6gbs
5QUIfm2Yk6YhuhHBIqaXOxwhoqquVNv1NLMJa7C2HRcDQJ9WgBEzdNbZMWbJSw/QkO9sfa2a0atz
6MOCnN8EM6EJCnRJbh3KfJpUySgrsCyWqMu9TzmHQj92tNEficxZLpoDILmS3rdbSldT+z1FWRDH
aguN9jeepaDbEqwjc8Dz+VZrjNz8CNDIeFp/ynl40JCbKJiLjU0GYxaVcxzocRHQchMuU5kh8C3l
6ElvED4wIsBr2yGqo2ggB8JcIPrqd0k2Zy8TVF2HViJX8ggu6772kcTa5k2LnBuaMrRzOI2aizKl
RCUgaonYL+GDq87P8MU41eYcOv9Q0D8xqGcr9ipG/A6tyyf4vGh+FdCGXEoOFN8yWwyMuwFGgAdg
h5qAUu+6/cM95MY+dAMaHbsq2/jXNcVeeoVKMpHJoLwd1ZLyjKBDEwKblH0QFaNTBkSo6XGpWqLK
JhmoUZ4vmjNf3FD8aCTPIQEeLHi6n92ZatybbCBt+AIJRhWc9XhVJPpG8DOUQjfU6t2Zx0SkvSh3
oI+kcdf0o0Gq80Me6ge5vRU2wgQmgTJhvehvPFudOL86k2VuJFmvMvfAJ4eaO/8Mxy8G7RAhMRBi
/iHxkT5VQEK2MaBUskjF9HkrSOgRkGDzupWWEmrw0pE+QG0yOmf/4RZ4fj++N++v8NA3HNK1UfUj
1usAkXqU3lTkcVnMfyzthSU26SoDeVq4Arn1HXHxvdNd+mZrnak7lp9itR4jY5B2CatiiFVqE0zi
HsvuCdVwodmJWzlc3L6EMs5kefEhTF+0Wyvng7ySHBCLoDCUHyjnVq64xnKDLGBx6DdYK0OWgbGg
Z4fHhDF2AOZ0oyrLkt9734BZNGbmQBIMo8bam16TD5nqjLJVaKnGsY6ymWNPgLJEwdWvP7ndNAU2
sbiZp8d3sxtMiaiHSUDYwfBuFDbs9U1Ai1zDB/1CcyawoiyIRP/AicY/yU8TmR3gtDz+JGO8LLOr
XzqprY2i6NUZ+uePOkMGbo6SdoptKYsS2bkHRRDAS9vBzemH//rHnj5ANlh0CbA7mcUCmsrZeUfP
MoXY3f5dv3NOwncoG7HU5cQfQco2l8cBxN06ESB56t8gviAYAJrXLyi8Wyza59oQDqSWCK6fSTqo
ztNYm1wNCjCoRn7CvkmUgckMhnW7b4MNy7S/CISvZ5KsyYVd3Vy8fVaE3xnALMIYndJqGthd3Ikt
MfwP02NYJ02Fr0FhRvi5IcL9tcjqT3EsVDc3jp6Xxcu337CM5vAFQD2YtiCpqhOiZfm6gHq+dfC1
z3kVUkJZuO8+msdjVmu1yhGxrqLzWmntZnMggfwIAfMCvZbyojzGe5Ayo7tRIh1hl3KGUWt0Iu6p
flMO2n5L58hsPjg6M98JFVmmRJ6wBsJlyzUQhE4zE3Whbzv60ctn0AoXAW6mKjgJS+j6skFL8+F0
mjKkNIS8QkWVvCdtA/pPQGL4u+7aB5BI45zJoHsiWUZ8xaz9Vq4xV9jYkbcl4Abk2LVB0/R32+1e
JkXXsrPm3mJd12Nsm6nchz2ygED+AQLj5JVTZHGajHVG5OPv7pYa7k5pFNshTMQIn+kQnhyYR5rO
fLrK0GfUhSH+eSWfBm6+WNfAAIn3ZT6zKgfc7mw8FrO5lNMM3ouyArIbgo9wut4fLGoxjiNGvpuo
ZFbShoWRBaVQAfk8s2dR0PdbOE6ZSWi8IBNaiC3uVoYRw5gNPKWssMiWFuNe54Y+XR8PITKs8hkm
ZtHG21zi59BurWRdSRtUKIsfUf9iK4hwAwDACn/RnZD3wqHH38rHejIioO6iu9wqmti+1IZigYs9
H1E3zxze9k911yB8EXgfNTcGfOhKT3mEwq/pmdKgpzFQk9u2V6ZUvXr9KUAv1cTqH2GIp+yGctXU
P7+Qd7XQ0Al5CmfiicpbEVJ4MAt0qd7c/0jO30jn4gjDHsi1T0YjO1Y3ePYwi62R/wq5BegKuosP
kmvsrF2W8gE5TgHc+oIPNhY46a8Sbk3d2N/RLxLJnl2hK8mYrLXp5C2YsHcFkUoCsr3lFJ00K8nK
+CN07D+C6eB9XH94Aa7dNQuh/H1mY2OdHKvt4jGDkI9vXI7S+kAxOHKVamuM6WL+KfRfWEFkUbRw
fRfA+FKpRlc2dUz/+g94uBsukP5PAcbzGIgFaVxyhsiGhLSaRxm0FukIa15/7ZgLjGLOv2C31l/b
nBwDHD+T65aQX3RzUJMMsdQZh8Xg9PtPY+84U1JsOrLmNXkXufwV638uFcfBgwvF43rHU8b+22xV
Z9MTekuJ27lK5qZdfGiqHboH/e9kW4BCVxngKUAwP/TmFpk2RUCJAyit8BOJIPt7m9+oIilDM0uT
IjJiqQF0P9/EoC+lO9K1KL97rUibg7Cqpi6A7NRMr+v40iKbdpNT4rAQvzgygADNgupqnllLssBP
EhW2JgI9KX57aohPFN2xQ0Dlzthab9IYCwcYc8rqVMLM0rHV4KZ541AMof4tW3/srHXA0eV6DPE9
1VubCVG00dFaqwZ292VFu/f/1zvpE7+2RK8RgLHUnITJMjZFMv2kuHQ847itiNr+8cvkEZnBMg72
y1kHDo9wWUPGQ6tUoJmPdMJS8I7R9p8qAxXXBirIcbDDvFSGSPXitEJIeDlAZIMWhf9QVQ3T/oPm
3zvXlBpELwbGd2Coo0PoKobooI5Yz+3koKI2i5wIahSL194QIwX23rKLakZZT1hY1ArUg2KAwCQa
07Sslz17iigd5Ai8YSSevCGZaEoUHxjPfx5hRgH/HcEgLBJmWvoEA5UkY4JTkjHXYn7jwbe1ho8a
q8H4XXb5qIgg9oyaV2trQo0bGazB9/52wBzh9ygMoIQWhAI9pWzkXKUOa8Jl5fYdSzyLybNRX7sd
i/V8t2JDZhT6N1bQzWXI5L4hh34XbDydrYx5ADss5eh+erfC0WctUVUtWLVtS0C2F4cjiAloV5qC
Jukjv1u+GskYVtf0XhD/ztN6ZFkYy+W2oLD/h1uF4IlhxcMrk1AxWJMyb/hzGschB0rrr6AhvkEj
DmmH/JufwTwZa5F8zGR6ZvrMut4i+rlXpFsi/fFkynRaNvmNM8OmdO3zQvLqUIuQzURV5wx31PRn
chUSeZQyk7D5sxgH6wgV1SfGuAu7zpVBUKU250aFvBqh2+as+379LLH00CrxYtDAc6S7PWZ+eJbp
3sAEFwHuXRWwixn8jbDd7zd4ylh9x3Mx2fknvane6T5jmXosf8PVT3iUWX/p4jY2/0uC/0TBvmz/
uUs5upXzvMioWk8CzGt66oLXrydxJkGlq6lbaK0ckpFNENZARiUScoNV4y8AhjEEJg53HZzX5L2A
5OzNKYoRVmGzZQ5SNDt/aGNP6NiK98emU7O4vEsYbRDHYtPW9KMyw91I4rEwcYr0ZymaCzghGhz5
iM6UsmuFjrA8zpukqREByN+uc1CW24WvG9AY1pBX+2MERSo0JVeu4SI0ciFvR5w6PnMW3dHJuRJv
Rwg8XRD6eno6R6K1CebPIRXE4rIQD1lAqsYTpLb9dE2geCry+2ZE2U9BA59uH87kWRsduxrCv11i
EkdwD6nweq/CjOWjGRFB3xF274SMlMmAU4ZIt9HYjhCAD7aMRfK6y87cXVvdxNGRpv2FsHbgtXCI
0iU6A5js2OVuWuGR1YtczN/peWsSj6yLgJ8MZ1IHtBDuETFr20YKkOyVk8LSbIQHqujTM2vTVJOu
AMuL9exI4QrQIyUoLCe4XkEgTA8odGds63SGTpnEquPX1HB6WPr8W/VYQ75Ibk8KswnYWNAOAuEj
CBmV+AraVdvUlO0YjorYfCEXwJkUeiI4wG8GRgcEaXEOcs6EY8wNUcPgkopAwJmpjOPQy3rZ8WPy
lEaauQf9O4fL/xh9UMQ0voA8KVwShmTiuGb2dmf7ZsvNaow8Ssev2wzr5Z0CcMATSERWCKhIZwpM
jeCkI4rhwDTjRC21jYABuJl2VKmOpwlGOliOnjUBHGvwvQbWtai0hzwEfibFvWHB8iwKMk5hLEjs
ApLgLBnHzb7zGotXAOhFVhFbCYjB/l/hTTYLc7RJKT2J8499elv4OH9sDszhXNeJbPwQXgWspG9C
e+WHUOQiL5QLfcEhiYVzBXeee74sBf3XQhY+Z6cp/f3Fq8Gcsjao9t+4EGpF+DTP7YzJRpp4stL4
yoNQ4QXH5DlrHVt5DiS0rCU7n/HRPKaCzIwf46L/zrxCamp+TQjIv1JZldLY9+GZM3pjK0pT9Sex
PZpLvyPv4yIGnW+QHUOqcNCxytWMoEc434JhlMJNhq910s6VbuqO/aKYXla6tyymXjvUEsT5edh9
wNiytf6/VaAZ9F3Ag3S1KgT05f+Az6Ie9WHyh8oD3ECEL81flhEBYb1Y2ZvVf50vol3ZFuumGAXG
LPdnKFegoFvp82XqxxjRdsNeK3JTaM2rpUAMfcXpeVhFAXCUc9SF5VTPMrOivlHMIm7SozKN1lvR
sJTwFalxvM74TQavO3A8JPALp3BVb1Ko7hhVt14ZbChqB6kK0b/ULTrHLh5DVtSRq7/QGTviWza/
njX5dpn1uP05ONrDOckqbLmMGm9/TBpiofZlXTfEqkR3e5gdz2I/RbNGLjWEjQ5WxiyesobGApjj
DhqmWhuhZYcjo0I6ijdN4dWXGgJ4m9qMM+JgRPiauKPb+RVn3KMB4dQyAhPUgt9n9yeMMWZ9MHhj
fQmzuq0bXq9r99ARYzyOY4caJePs5Zz5Po/UEtzLd/kbVXN+HwnxQNkgd5632yVP3NHpubGA6oMW
U74QOLniK7BM/L/q8Sxawv6XmQyhw89WrXgCLXphWORvHepAEyKGa9j10FXBrtYyW5KpInl+1ocm
zYS7MMv1u005ZEyXxDFPPE5eLZPK/QaLCw5Np6wPBHV4ZwOQjzNCMiRE0xX7wFpmfAj5mAt3kE/J
ufh+tARCl8kB3khAkXiW915zZjgze/ceapWGRBkTeYzt7YbkysE09UOzhpMkdJuHg+7iWOSKlvkj
sN+/tUgSumRDfMMZRbUVYRoXAyOydMYL0TS9dqHDcSfVeqwgpvAdME8WeKyw7DL8QyYQc3Dlqx2O
wortiktO1Y7tYIEoUE0BMbLluPO8STR0u4Lpb+6grOKeWWGjIlPPIQv0/NccJ0UFLI8nTEDhRgzv
LaPBEWZMc+0uHxe6PkSvSoArQMveKzMMF+0hlzZ9COuJVOYdoPb+D9gg0gdEZmbNNNjGdy837+Cx
+2l0hjjxcuF6TKSP+AITwOy0eiiSrDObUq3lEyO3pq7uyBWBeSVTmwgAgdwwCTeN1GQXkjhGHwnr
BxpR/a4Ha54Q+CD3i08sS3DnDITiPt59GwwiF3czN1NT1+UPwZiRProFEh29jbOBko2n8bepdeQZ
Cuhdp7jRl9b+Q1r26Tr2IhaPHmYO1XeNsVpeDntU4z5slDYicRLZk/qVD5lIxIOi11tY40AqZTpP
DGYZFcAyd/hjwHwv5jr4WtV7qcJ4LsFg3t2G03eCkP4ng13a/48DmLnFX6yr5uRfwoQkep3AvWuX
rvJ8t4O6dcn83VOZYNR0Ts3ETjMGAq6RITs/MRq6wxpGglZqdbm+8b35SgmYileYL2w4AgweF7A9
i4RCv+8jQ3xm0cw6sxOGrxZVIlN9yF4OJBnCbuUt2ewUrs3GvHh7YBPRzcgwcfOAeUFQhQ/D3Mtm
sdSgISzilbihJOw1LE2j6/zxQ4ifyu3wT/nrtsDs/C8e3m7rrH7kFBWJZ6ydgib62zKzapMqvrVa
vJ/QawLNi29E3FlpncujDPEqOjwu/6TN5EdR+SDLIwrWiJh35EpAlxCpfppc42Mlx3Z6icFuNwyG
aQTfcfPWBt0sQ170SfF4hUDyX8Eq5sm70U8K7guWHqB8Lo7JY2ZCDITvRONJ1WBm0kbIYn73su1w
ImAbiPpeUcqX2LkeAGKhxb4cL1UTBwjZn3m06bgA5smbKCBvoKNG4YMGGZoRmx1YWxcXdZMGdtsc
IxflTWBtURq49j9qliUH1VF5J9qAAU7vaEggQ81LW0abBnvc2U67HHDSDBa+PwK+lVKUfiw4RvpA
7DH3c7eIK+3ezYrBUVRrKxUdds1EMvJHw0DlZEytq4qmf8z97C1bjZMABGYgyjFHkY7JByAWe+GN
GiNEL9noFcPC9DPCqN+7oRX6zdxeeQ9Uz34MSsj/k0iAFh+peRp1/wnuGEf4BgdfHWErpnWrVEKR
nQxDmM0HB8QYIooW084u9cpvV+sEhs7d37gTDkfdwj8CHrg0VV1zXMGu4QDFj6G+C+6jCk2g24WX
aiTmhkKdDM1QqlraEuRXBKoxGtEeyq9ClpsqT0aoMre/XTKz6UGfOssAK1Cwt2we9dfg7pn49bRa
SfktZZ6WfwqJfmMlrKrqvUVilNbZGD+0edkMD3xz2HhIucwXPs6DKPVNvuySyiH66UNAlRaiyK0i
wpuPy7EmGJcX9Tg6pg+48f3qX+0vPgWNJ5speTVLisqgOCWLd4pRb3M02EiL2g6CswLOBQ8F/77M
mQwY9AFWFvByyom7peDu1otcUuPK5Ss3JFuJKkA0LZgD8f9joWh67MaBR8In8YPyH3rXGwckYqpX
+9n9rXnyBIX+7TZ2163saohbPDmfC0nUU7d+7CvAgrNannWYeOV6q7bwH93l9P2iLKJuawXJo4CR
Q/Hm4NXgBz2+m2gFCXqP14GDOttgQTEWMec/vlOB2nJ1J90NHKQzqsZfMJ2Q5ST53hAY/E78VkIa
/oaFG8ZwtF0ENx9uVgYRQzlJZ/cHWxpAT5Dw32ZJuajnpkn2iewjCIB0bEra8+92s7Mar175Jg6b
I0S5vL9b7W39qnyL+21HYJHfSGUpPW9Qy2F922BxBVEWGigJPCD/Oe6J4dXZDYcAKYjzMW+g/T8y
t5P79fAQjAm609MllK6xoqywsXfNjof/avSf2UhoCzwZs7hqOCa1l0soP2mKP6GDX730pL5tYqaB
ug6bq7wOytdpP8poHnew3ICDmO/CZrIMbcbX+qOWxE74yTrsxC0sX+HgSRcywSCU/QfvtjBuuoUr
HKc+yJKG6a796dmalU578XD/QU2iHkRuebWEnJp+L2aUopB2KFCpsMDFjpf2DHfnKndNHkm+2mSR
IGKAf+dV9YwCJ1Gidx6IOGj0ZX8lili8SaInWvnRr1sFEPkSEPSsgUY2ReoV+gMfoUHdrLVUZuGY
SCwPsXzlpIb3QSr0mPMoJjjJizLC/tqGWr8s0N4MeVSFpA+/caZINSANMGo17IIs9eAPgxNy9ZB4
TcsTwqE7CBAFpa9kgdvSCX5DdVmsfSdTCGcn0UvXlnmfu9eEMlE3HDzwY6EW7w+TANGsMpvSfdM/
6NDD86cOpxWbSaakFK6rsGZXir1SJsulIESNJCKfZw6wZCCJ7vF03wYzs+xu00BPHrWaaQv4BrYO
Jx9q3vq0gpGZRSKjCZFiS8O3ZyP5Oa0uTpn1rr+d6v/bElib2lje4ym5sc5cS8zvXKPZFXF3f/c8
qHNm4Gwy4MigHCwHniptXR++XHoDpWcK6nmo9VcfKeQoudIFYiq1oB9rtUj8tFEr8lmJ2ZEs3bDa
BOrx9fxWRI6SNzSWp+b7BDjRF8gVyy5fLpmkemGPrhkxuy6HJAznTiXvFziet+yl0AcewDJnKMtk
2EhVUrrFv2nmwSnjJSW7A1Q2lATqbS4cAV4MlWkgEAHRsN9cmULvodBT2GEoKX969RIp3U70I1bS
tHwZzqP/jiwifJmbg3OidCXucM8cgo+OcimRGtAsUo4ePxGNCV+2C1h1yYdK7pfkvXQ+P2mHjhmd
hdgajnM8Sa5Gv+vBsN78oca7admECLkwsiJ5mDKO4FCi/LGabkSSG/S+B4ZvBAa9fzakTkwePfRm
qjmPWfDX4Ca/1FUrkYw7D3vciculM+OQPiepM2V0amMvcQfqhaaf2L0i0PEXo6bGQlDJV2TEtuuD
RU90kFgVxs58t0E1hUWYfzTplyQ1qT91epCatORMD7EN8Z4DZSrvAdwLf31xWC/S/Cgn9KrsOpS0
nL778B/tFXNWOaLzcjbbp7TP1RAXBUvnbAp3ypfziSRB7PgsrjNHt70c3Dnn8p7OuNdxt11YdU7G
WJACcAIPxNPuCuo1MWV/6t6AK+kfJy6MLieBtnn+D6FEPHyDQWXEyAY2BF6Ybi4xsy+458VFqPd0
2wzw7wD6I+4X5Z0btVV+o7VRnr33Npkp+NVzGJDlyO4GfR28IfGu/toN2AG0REcw3FTz/N3kv+WI
0YKU3XXUAcVmdwp8GuhN2i7qr2rSWPLtcsRewUL1ctppJB1lZwC8LcrauIMjqA1d5Z5n0GlyoPeQ
cMrFrdcYQU3vy1bEcMBnoartb/jM+tUajDM8gHwYoeB7b5MuwjxD6pR+27wmZgeNkeS/GCWTzlCR
oSG0+6CeIds3IsKyUw+C6H+eq0FYKdfYOZYRUWRsHZZpzxEQQe9YLdu3ivTpia8xQY0cgIE+hOJ3
mox0ao99IMxrDVufaFxIwHBCvj7SWqy7Pqjb1AnzXQ9Lu6AUnSD/cPrj1vQov+Y8AGWVfNOJRMsC
zTjUDmDKS1zGEtSZGc1046Jw+ZgxKhBu+s4gI4H6LGqcHgXFUknMV9/Zs1YwxEocDqG4pevY4/Xg
ClaGRZdFi17HwucvjvDCO7wzEshgxndCFxwBrKGuW1nPdvCzu4+4Wz9IEJiGYOREVFZc467f/wLv
4sT2rPr/UG9FSWOFWVha3tgO7d73OvZ/991OSrXGF4ottnxREM5wObarHxSgbGCat1Y+2RSlFHBY
aJnkJEB9jBvQFsLk+FTV0itBcVzvJpTTyHqkShTUfGqUvQ7GliOYA4NRXgr0+7u+Yabu5rj3WQho
w7PXNGKoJu6jdvZaeIoEB4Ti5FoOXADsxCbi/dcjTBWs80k7wkb8s9jM76IORtLiuUpglEaw7W5z
w7y0ne/NWgi/HTRMrxZy4+4Kvyg3G8D7EL89HDSOmBx6U8YMYue//z7wMi1tUBS56Phl4wbndGG8
G6QzG2hO9TfsfNHdQMY64EhTOOCuB5bW9IzoE3ahSQ+uXKJK9kyVHH42Vqy749+AkiOANFLDQTeU
lAL8ZL6kfIJV42jiGwdi4km2vhS4lV3wxIYegs8PYhLEwhIH01w4nacVz0n2KkhaTHbNQhYjkSM5
tS+KboTC5lrkFoWqSX2qPHZttKJKCm11+UUYLfpwdc+a6xPK5zq91jzQ8azHWMupylvNAvjWFeWO
L4eqPdzaf6quGrntRS4eH9tF5N1pB8LZqNryQtM8BkTKUD04YKtXzO87VcD3wTJzr5cKySFZkjPR
mnKp1Qj/1Xs1wyRXqH8EdU607zvZi3TrlP5gH42GaDOmo32LG+i1x+JRH5IYOcBp/oYIKLEJQgo7
0hGvGncp37Qxa/KlstXRC6XfmH6W6QCCGXyik729z9HoauRilL6x6VQxqXYStlwHoG8/Wf7ppKW5
VLb05Uxk2Rp7ThFUKVUswVxdCZekIm36fFGuCpQ63QSlZd37JC4mD5sjxTl8acrt75HLTcfyjxpE
WRVv2s5dchT8lawUM1ua8gnROq/mSTFk0rjZjcDPUVYkuTe5qx2DTLAeZahpIJYyh+g3kTF+LYjK
iHWiQAL4zagNpjF86+zQvhYwnukHsMLXjgCqQBVGVe5rhufnT5VffR05pSrEfubyWcUyB4x1TTLN
OjO8OrjT4R4CTF8InBge2+Y5MaT1Fio2EIpA3yQ1VcvIl0IujBGUF6IfCOvsqyh4BRaNMb8Clyth
DVRyo0lA+jPCSjLgh/HLzyTZD3h4FGArGZCp5OKr6Fgz5F+TEnMgQlhjQGuxdLipn+YC3RyPGcMU
htJOa1Bef91D4P0KaQS0u2282IB0avfltKeGWhDD1/T8wvSzmcQh5LfK/pF3vH7Pr7w2kPZ2LhX6
RkLoUMl4kQbFFl3r9mYbFU7I6K2421rrYd9AbDie443HtWTQCsEMORPDgWugDpdsUe92FP/EBvvP
UfRbZhjuyLbMDD0JYjyt4luZxKbbrGLi02bQaKEds97XZNFlGZ4k4FPDvzusmeuUumkNELyROBex
8sKfRRXn7LyXAdV/Cv9Yrqwt1q6skDP0HQ0oDcEvFYbjeXL3QbGxYcoH1/1yrJ0vAASalC0kO0yn
YurerAFU6EkxBrxLTTQ7gopYHIjKGzBk8QKf9g8sXlRzZKN3ECshTrTtQTOzX78dYouwwuLMFluc
5DurZIbBNnxEc23wNKa4y83hSNy2QR1lWVW8SLlu1+76FI2OY9LfPkJuHOMv8/9OzU11Q30zO7SQ
1A3guXjTP86Js2cJK0geFWj18qaR7by126yQgzWvhchn0hWtUtrdr/D1xy0k3DtBXKA11x2abik+
4+gX/BZUCGSihwlXssPMeD3PeyQnnCDv4fB4L35jeV4RsLp2k7efG2aZYZim0Ss6wlNBfsQ+pzc6
6TJj6hNw+2u+WKNVcNRHdgFfCOBDJa3xqyrE0v21vxBeiqfAlb/NhOZAhtinl3TyGbj1enAM9q4L
UvDdv78KnUqLDQnlD6E5Sr/jXeuCQXr2Qa2GSJ4aUHttN3W1J++5jD/HlykqlFFyavj/CUnglybH
4rEFxwEok4h8z+xzIS43BdRk4XKY4GMsLun3ocVCp78FSwkMP7XUxGkaGGSEs7lOIRtjinVQVer9
LJxJInZTOJuqyzqzspWRBNm8Ts6+8pRVNVZaBnjsRg6E34qNvci30538MwIGiIWJdIQZNuxK0yoC
cNF44BotGpFsu4ao4vG0PhFY6cHUdlED+Q/XQPXB6Vx3HUUhhwe7IbrdhxUcrk89IIM+ickmMkuT
RzpLli8HuzOzzK94heAKGRdZRa9l7J8J92d7PHUPkI5L8tAK1QX8ZVCgkXiYl4gKCi6QSrYdQ8M0
PVNw01t6uFAFuF9sQk46Ch3J6mq4fr3kVMp8z6DigTgz93tiu/KsYRBkLJDNWMAi6JxVRrITzZ6v
j6kKGSBQkWkzOf3gBqeyAqr0jIOO7VRT/4kXjzvg3VOCef9V+5zFafQU+pmX9dPNxlgpecqBHEI2
jrKUifoA8ga0mALC0U5b2FEf2n7W0hKExCWof5PJZM1C6kpPJC3dToDvfgH6LWaktAdIkfxe4XIV
4cETqoJgPrTiYSk4JymQQjauXk40/AKztiKWlF/+Bql5MPY5FpA90/+Gb7wO6hsbicJLGnapgpPE
db0soZE1fJx935eJmjuxwYOaidBm+a6RKyW/peNFHXeEoVQSlQBO48cGyKG0K6OYiVQcjBUHvDZ6
4VzdCJJR61E6xiaOtYDX03dkGYYf1ap8GEVFeADZY4FNHe3P5DwGQybMVtiEK1y3CYAdQRYZ/eVc
OqMPLaYwJoMEkachwbau0QbOnzCLT+8KuMQF2oR4CO4Pber5HE940yRRx9tXLXyuRqWjvvVBSFh0
WArxAga3ZCV/Z9FNVhRmmQ4j4ZZDLmu1l40zMB5lOoVMwAT/iWMmgHt5aDKN+tZVntqvlRWEC0Zg
Oy5jYwJ56DfXcrtfuWyCFXGzNjCFIfeEMhrmYnu6PCsa00/9CVLnXm6VsCyrkd3l198w3M0wuopn
P8JGKem5AYIjsI1rRe+V2Tw2ldEmRj/Vv3ONnF8K72xCJTyutwy3mZYJp1Qd3+1XZDVh1Mw0JRjA
K2PlTop+QwJ8E4d8Fl5CIc+ocTrirladrcLZVWOWBHbD1mHb4xqsREsrOQ8jlSKc7uHbxDFo3PHN
I+1wQY2sKdRyERVTDmfExV8T97dFozcuKx4xqEh/Jn+B4lDhrId0iCYOSEcv/P4JfGqO/hDysvK6
JFMLz0yWzvF0GukqEI+nwCKzNGCUhFEOOpnHF3oEjZ0LkzQuRo9TxdnDamrQppJWvO/C/cLCVROa
vXrMlLewLro9fea4Fhr2EjVwFHRV2WT/p4HIMhoYc+64YseQ9Kf64hOm0Q+bg39h368Oqw2PE3nq
0sXZybaE5jvY2TPlW6gzZ+qZku2ltIKc/nEnWmtob+jjC4sSXmkvaehK97ZHHI7uYJoBqwCRojGy
SH94hmTg75HqVFvBN7pkwNSETKiAERpp0GcXIO46RjxrH6xgiJoRrZ3TCwVMNAAaU7UyZCuHhaNv
hgxWcYWlSrRcFOhaIZO+MumlgoCKAknzPkMoc4+tklFQaN45rkyltiLnw4K/Tl9kwVDc44Ejfyt/
K30W1IsybI9DZkZTDUAma4TJkLA5iJ8hcmssY7zbLZVWaIShrIf4JnNmQE3ycA9WFeLpOpiv8HJK
HqXBXyBNlFO74+8VHMnIyo9H9/UNjXOvS9HhQkSJymo1Y+0n7Z4kflbtfs/EeWw/QQHJbCEJNR8d
tI1oGKw8LkVkFMX+VD/cKI4aRHwP77k2Q3eMVHgo06nBVYVlHOii+3V2ydUYMKnkZaS4gAP9wsI3
BI4ZZL5Y9p9GsrF97xG5MNL0gcqux4hACNI5L5Q9D6TCmQaIzAydE9DX6Cs481Rf7WejmRtVbIYB
w2Eox79lGqJjU824+63kZt+QH33zTfiDWJ71Bey/tvGMHrf6CbLTnD9ka4ZcK9KvSAJS6JXGUJsM
NlnREuCDH5hPSb6H/ppSSboGPaetIgUrss9T7B/CfZtFzJSObMjNgnAcjSy9YFYuVWBMQE/wiAU8
tfD4Y39LjjtN+9y8uM9qb4eHazXI3Nu63lczc62e/gcQ/eUu24nX3WvT+RD2tHJ/Xx/LhtChRtHJ
DV6FBfL+TRNdQhfHYUHA6jL/NDRB9zwZD7hNr441eRVrnbOOFD3pl3x7rNw6bnUskE2hL+jHX4K1
tNm8Zuo2qwo1ZJEym8lPAOD1xStoX73XLTvBtTlJhzsX/xfSo+JsNhQ9Pa0hWmkYyOtb49N6qr+B
Em3fzAYFv213G39M1q1qobsCyeARf1Sv3RhEGpJckEVuBzJGC6z2OiAG1t9FoEIw+l2EFytmar5G
G8QMxFELxdWp2YA3sCVKnAlL1ow8PQVneeg+M7RNNwUpbOSVkLKisP1aw2XRfxIqf9OpNal8cOzT
rqfsHgA4NGP+TykX/r3LWVFW6xLaKP/7hJ4TI67pVDcsDTjpXLtNCay9ygPb/1JZpcjXzymAtTYj
CpJMYlq7FZyYTDei72EPmNMaCFLhXNuGKVBVY2fyq4sYASMlkC1Ds/1jf/UUs9bY/NP7PfPfKZ4S
s2zTfPYDTGZWkrTsHVFEOSZLcmC8yc8ibkC2l1zbBVsuEZqnxw/wn303tQmI/6yVeE1DO1An0At0
F+kT/vpQN3aS3tyEz1rdEhFyoCGewJf/mSS/1Kb4Ps9VJlLKtYTwATjJavsPOHgbfUTL9I6qazL8
tA6txTQzg3EHoRe3YLN2RfLp33GJZ3aLO7v9PRD1sZmKjhVo7GHDtCkKbeEeLvCnO3hCqfxV9mFI
86sht3Qo/fhFoXoEasECpxGtjJzfMovENd2p879q5vNA+C18azZxtEyQP8Cyg2t1nruuT3r/iRd1
yPC3wo9GdBvR8qpjIiW5gIDrj8unXz97x4LXVtJYd9oz6YfH4Oi+nICMY8Y9XhZFu5RbLAsXUiOS
TixfN8LnKEoCkj04On9DYre93d8tCe3Lq0eVsH2JIXjmPl897CuwpjfKJjADDq4AKlmMEudvMWIp
Dzh29+gQ2tT9TBlmQk8+CtpwEc64AJY9fiwYrO4/jWobOp8FNCbZY5h6/ZI9tXweBd7I1OPkunrX
h7ClQOBM4uCTHzgquKvNeIY1M9gWSnJecJTf6QTYXuh4dhC4/DQkdOXXZQFED2D/HO0O3gXegCMt
jnjz/8ncl1s5qWxtBs/2NIkwrdgIEd7vDTv6TsUW+H4rx+HynByBpXX+o3v0CFczRL/b38KJvvsn
XDNoj6S98qGejsRWzWqVdchdX1TkE7ZUFlq5J3YXiwIXzdxi4U8gVWWg2IEnAI8Rf0gKatx7t0lL
z7VFU0TgQHUwxy1Ucgp/z0pypQ1D+cJyqD1puScTiNdJfnSaGXYgUNU+FObWrTr3wUMclJPOXDfB
TcjeE1adkA9bNVN9BW1RNnE2swMegx1xZiUtPIfpguphch3kGbrVaDo1gdHyRUj+QC9t1mjhL+K1
Ep5emV8pCLqaCIq1mVVpKJzeS8adInLEQubZshDFspYrSBbNpnFPGvZDDE6sZQ6KOJYXEA78BhSE
epzwYi6gzFwjJcIsGDdM12SnxnT5vDxD1G8pJ4KgPGgiiM3oW/Ull9i+QTIXhY0ugQWrBTFPSDzk
HpEub1IGO20gleCz+Asq1OXSbEMctINhZVdphgTXcMvaCoWrHFCR1231/aLLrYsODhcERh1lKaA0
TOjm4PeJDoO1Jag0l/IWcI6h/usdVg3wGpYcV5pL2Ta/fAW9dfpAidq7e9UWdx1DyoZq1Dcb9Oul
TLGPX9YtAnCxTwORmaPrLZ288gN+3huj1pmDmwFEt3F60OgNw9HL3U64voHn9OiDAhrr408AG0Jv
zrPoTZAadXE4U3iZziUQFNJCUdI9dWzM2DOapGUtt9gegrX8sXzSlHTWB74i4ZlB4X8Kn5DPdQlu
RXhTEvwIJuP7dVVsLAic0/YBTxPbTAwZR+kppwxmwzGhFI5FIWRAUntN/kULdg9E5aSM+/k1mbL0
Wv45kWtQ2APlVwBOyQr50OgPjyP1z754ttPJe/1RksTc55OFyqv2NJaw29Itk6LV6kdSPDhAPHpS
Yn2I3/0c/SMOwI6fAoh2SVQkgSjW7u1c0WBR1v3KPzFsUblErIcy5NvNadQVWlt9FphXAPIkBh2Q
drzk6/704CJ5iyyikfDJEcMorwh5NJZtyEp+IqU3R6WcckOSj5uUnjqsSKumOX3qqkUneW7V9zQ9
U61/o0d8q3qzkoVMtKtVa2gTVAg7Ud3WA8v3IGCB0NbmF0UyRh/jT7PNXiFLjuzdg3MJgxUFKdAl
e2l0by2BNrHHoS8F4uMPB8RkX2XIqogstBzstqT6uvr3ORNconC2e//6bhv+q8aCpubQHFiqv9hU
fo7Inxta9Tb85+qa6ngymbFIGg+loWpCly/P5L+j/xUCejJhSQC0sIFOT/4I7Qudyr+7T9UZ8kJx
l3KIW39ThNlLqPjJtNmzdYb6VPyGfXE9oXS83AiDvR1m1qv651nz6nUOZ8okTcOu6srFslM2l/D9
XM5OHanwh6QFj15jmom1g/0v/Q1G/S44wYjpuSDlDmmzx6BQIPY4PlZb9yzNBoRXRTdmYcYDoEby
clbCAq+dLPWlZZqoe/vyhZ8s5vi1x4vXGO9gKNMT5HhKRqAze7oMqGQvs2VPjii5qJ/YwrsuXv7A
2wEjlrJ5ZMgogjl4BQf/4iWL6TlH0EMBQ3juU+jC3wbUgvTiXWgKCy9HbOk/QLJTZsMAGadgfLkD
eMuNKA4h+cDrTMQB/u27F6FHEcV/8OhoSurDfLgER2/TiD9514Y8hkBtHk8+2E+VgbPg5KZln9zd
O+oR/rLPR6FcngwiRU+7e5B87yXAi+KSBF9eOlDbjmN5UbdeMUfqlrKRG7YC0CW8jRA4jGHAkIvB
xpBIPwzbVdWZGEDsfiaxQ/leYBft6Xu5dnNDNJccAB+kNuyc/MYW5XzVJKgcX77K3SpDqSjtN4Is
TDFDQEpd+H5vgWsbv6uNtbshEwXlCC/8KKdnf9MsPe2J7/zvi3gO0QQnK5EfsA0fmjM2VKQLNEob
EkwJWJZuUD4c9n3FSB6JjhtUeafBc7jdklSHxUqs9QsM8HafTCxPWb3OGTGc1DFuWmqhZxI4ieH1
TYevRaymSkfhTPoy/YU2+EGbHA7TcmaoztnNDycRdrXpwAF/CKIqcocDYXVoZcDISv+Ss3x94eqz
+Ixcgmb2w49QHWMK/BhEorIUcx8XIQHM09h6nkGzbRLmlnZw4AEc4xC4btireEzjUfl4JmgkZh3t
U+3MIJIiXZ5vty92vj+b+d2OEzMYKr26hqzvz0Ts2m5y9inbPzqk7E5btB3kgdseBgD58PpUMVJk
nyMYgJu+YjkUuI4BSdgLLyQbkSh39fpery9mnpXj1/EoQIWTRpWtIFw7f45gTy3JQtAu588GRbLX
go0/lVpNoJl3wAqYqPB7z8hrmjg6QNYfQK2lr1O5bUTfVsw3l47op46x3w42ePfdYpLHiXYbxsND
8MHC+s06ooPwOW635LYkRlD4HAPWOPXW+jVS7KqaEGn857iNQFBaqrdDPjhCVfBET+q+oxjgj1qe
jwKCCod0gmtNR/n4C0YRHvVt4iStt2iBS5y4yl7egUA1IJQ5Pa4iUM9agGKyjXX+pM1l/AUw36oq
hd73l9xrBrkcNvPd6WFSDS8tUbOm1lE5v/C4PtWvUtvVKaB+gv/BciSXrnN41FFNyVrhoheD5Q2F
EghyhCAw2LOsKZBoJCchmRpc6agcQmJsFHwCx1xk7FYgOO+Qz5CB9xuOYylhtqchNoug3Se8JugS
xTy+WFZir/WMP0DCETaEROV0V+t789u9EWo4emz1bs4YOQ6DcIYYQZr+67yMNVLioyJlrilY3kFc
5mjD6t/alrwTc2+FNMtGviCzgJ5irEBNg+OOQRgQSHUuck5WXpPNw+HoldXiBKAg26ugrOylwqLK
G9VVsYcSkW+AciaTzK54/GfcTAhi+d6BsfECpMFXTwvPoMzk4hgZXCRE99Ke4aIzDmgHa9EHWo7k
A2dcLUJjXUx2ucrLnxvsgRjsHUgPKLnugFQK4lDjqa4nYkpyIYYevSXCXGeMQOMieHh504/QHy9D
8zYG3yTzGX9OS7fFcUOhPTJbpK+qARJ5YdSU09kPzKAbT+umtHHuoytzEeyQ7cUaw0EzSUjqoUfL
ZJUNsn22fDWvndstMmPeAFivZ5hDFoG/f98bo9tBSlQEcoVB2R83gAadCmUGs00S6Hgg0twk2sz+
l7bYtI4BlTAqdrj02Pz2DToMDQAjHNbW02e4ZY/t76P1Th6apZupLJEHXtSwTjczKtPWpkASqwm7
3suVcZRKeoJu2NLePtWeURQpayNjxpQ0A+v4VZ7wErY6+WDOz6rForH7Mnaj1sk4MVzeAKsWru5H
C6Myezw02Khu2Kd8+XZlxsX3mssB/UU+EM9FL//C/eoHiFD3b/OwezrPVikq/kyo8u1v6c9mQd/2
d62j5DdH4x1PIQUKkSomnagBaC9OaUebEQ1lNC1GALzMRaiCcbZv6ygF0HcokIxxIoaVedC3vo5Q
fe9G9mW4Wt7H+NGcH7bHlJFM8IL8uhrJ0NGE8ZG/pGmbV+fF2JdPLnBDaiXBPzUy1AVbCWKa022p
cyWbKJ6bOF0AkiPIZL2ZmA98I40vhkrXHw5k6ccIe4mE9g9f5jpxpkXkc2q701/Ilh4MemiUnLUM
IHrQB3SJaiBo3erQrM4nBnzks+CCNQmlMjXSXfpYRRV1lEgsMRsVKo/6r0L5ly9VW4dx+ofGWUMO
1+CVpCfVGFM0a7WyG9VAJge6jt9j/uU9xCvagO5thzwWU/TIgNwuT0PgMSYlpJN9Wz77oJhY+XA8
7eL8p6t2t63lcF2DSu1h7UXNdbwFwm+aMCqS9qNG5c6Bg2l09jUyFEytnJ9rnLdXWoOT2mPW9HZ/
e3s5+4AK270pMT+b3Tu9IlbjaPTAxi4hftWAriFgyTcIvULb8/dYB1Gz6igSBLKUDgu8IuARq1U8
gyH3e2SfDl/CY1PfuZpfwBMJd4PHphH99gVx/OQIWrV+hdwAqvbkOWO5Ml8FuDof7ul1UjVV9Qq9
ewB1l0h6TJhlCeADXxSIw9mkE4ItXXY9HiASjaQyZeCz9qvMq2bCW/FY/1FnmPXbVKu7/62tlWDT
KUAzNjgqXFX3TpsqXvu36OhK0EkRqbWAMTXtv7kQjY8Ffawdi1JlXtD6bRNX/hLHBHnGavjoflSu
iobNTBiAWcJYMn80UBH5hHkaUmcCYMtdRWt8jACA0W7Wvzh2oTDUXKlFA4p2eiNGliJuAVSxoeHZ
zvze/7gmwNdbYkZVRauz2JbcAblNsmeMXCmHhUQRjMVZ5cnXXQ83hmszlP7xC8rgQstpCQCR4XTU
pRTSbxcS5pOdDT4Pyc4+GYdCDQh8fqFzFhie1duOdKuyc4eQyklBTrFoMFJWWpWZH+28qlHSkcyo
W77tVC2CjXjGYME01ijG/ij8KadrvD6qW4A0t30w6PgW0WwrQspiz+uzDMtN+bsQwaBg1w87ukHC
8M2jJlMQ0eldg3QU1w+PR/4AP2gOA9Ez36vmSi/yYpdb9flMiaLvya6eG65An9YwPxET7SD9XdeF
ptzBpLx5WIMltjzmKkLWeRqur7GVVVlDRTzilydGH6DSLborGyksh0d/38H78aURM937L0zrZ/br
a58B24xZusouE2CrI+HAeJhEzDTU6GziAhwGjywn/JG34v1ijJWi9IqJ54mLgApClbN6dvlNg/OZ
Zx7ApxzpMOd+0j9lOZ7/BKimVF3eax4Lm9kx78FbsRKfXYUPdYV3CrIRh/qwNfGMGRSGRKooT0/l
2E81s+8fyjaUnhI15xuRnPwR5J/5cmEHxhFbAJ/RLhYlu8UKjJsxClCykNutk4Y1Wm9c6/zUe3Rd
5lMtA0YVkMY6pIJFFMgbKWKiIuag1RDkOM2G3GJcoMPfyGGFcatYRiowt5iWcfW9S2OIUaI1qeK1
ZyK/tzW3F/wuDYe5MEbdaodlZB5uM5wmC8OIKKrzdn152ujPMOBvC0N2/oAbWtFDOaIVs0uLq5kj
v2FRktinEo9ZaTGMspoFulrB8jc79yr66V+M1Hp5vsWtgLfTME+ZDHaBI/DB9ceBWyyZaS4pa6V5
gPUv4xt9Ff3Vd3dsakPbKpCDXDAa/QtOQ+KSLTJs5uURuAS0iLaaLIcZ1tgiFXJUFqQDr4e7qYzU
br9AklroLP6MkD4motuWKpViRii8XmpnC7H+NHmcfyr4+jEnUe+drc/vpTuBezrGZLL73ij9HHfd
3Cw+uvMweglNIbMX/zpvyX0wEBpw3cG+sP1lXcVUCA2dPELgYQZk4dg3eWMlHwLBpC3d2K560Krh
EliAYxd3KkIdt01tfCrC12rSdwKzZuEmVsJ0HvbY1LncyrXbJ2BkHofDhsCV4C/MImQeuyYY93Ot
pkwxjB16wAWhN3eSOVB4LgetaRK5MhhCcBlEASPEUCAWbQn031pCMRoLzYT0bANi/22bUJn9pAGe
omc/N68JzIK9xV5S+ibYoWQEaOLsrzRPonm5Ix4XIDooLwm6NpHh7hfptldfhKXg7SXAdheLd69X
zVpbFG1uMbskmeu0LxwSh7AclEE76WqekhLEwq2cFFz0CY11EjWJ2SoJyOKzmMNxYBNghftGuw+x
QPYR0A97I2kA50kgW/QPzgt1jA9+qU75FcLSj7TvpJlPytmXVjhk0aP6Boa+SrLvmFDqrJyb4BdA
92Seq58GzRlsX4LzRbGZSNotVE9J/0fdGk/UWA18i7KLGo3hKjvexGe4OVZozC9g0GoYsG2aO4bv
26giKU+PIbOtIb/VF9tvFMua8kkdO4dExYC8ddre0ktB/e1fz1ri4D+tO1o5LoCorunBCI5xbUPo
PjhU3R9/kWxihM6qvPTPq8Qab1hiceXpA3ic+f5NPswc1m4J4wjJYwg5UMKWwr7ripgkTjcFm8lx
1pwnIhpeMSdPJOVYumuS4aq5Y2CZwPAsRquHn/gEwWY5jjUkG0vmqpaDhCtZ9Xr+sewb79+uNdjF
h+ac1+/XubzGXsWN1L+Avcg6b4pYAalq+u/09Nexq6CarmQNJKD6FZ/0y2IGXRW2XnabHSrbOPoP
zO6/kgPPBOOPeGVujgErtWkbBIRN0ZrdBgbWRZRuLE93oh+v8Whl3kQJCX1Gpzqk3TSojOjADxQy
ah8t+y/+D+BNA6hOtK+MasqhqDSi4btP8f2HA4s/HXtfWJxrfGbaKSd+uHaZP0MtErpR1qPzbFkR
VtlGwBjLbksrSdIIxTFdujrx8wrSnz1e7dvJCa/QrZj5htp7nrZ/B5+UKC3A8L9yPeQ7H19BCorf
00VFPoO89MyGctNcH5ZmEytXVcC9jHS9CfaAqbJGbsJM3XcRm1S3FrM9EPgelwoczzYA0yvEXrRj
k1dMZrTzcJSGqz8/Q8Ms9mgv90z/S9sofezm1gWudd4Qqtj/1YVILTXzHaQuOWg9FrwA2QG8kZ7w
NCya9GznOOEsT0akq/bcUkzdDzrLAJefs8h6O0Xjxf55EfIkMhJdb7Wpj5Ac6NQmJPVmQABcnurN
riHd+V2t3+AKp46dAmB8DiC0USlYUDGCjTgh+dB4ju71ZvK6A6NK5xxFgQ2LfsTyq+YMs0rRvul8
EpxqROhvWK/PnsnyhXGD8g4B6SpVwGtiqcZ2+R+wnms8466OS4DJTpIpbdK99Q+b93xwte4qaJbi
OL3tWSlaP04vUmtDkgesAC9maARb/bxkuYlCk8PzedntG1e4cGY9Ymxgx0wo236LQzsH2crH0Tdx
qLd7qXH2XPfWLKKf92VR79NTwyJApkfEvIMN5IqrUbWc1GfpGn1CoyTBm8ViNIK0Lt9MASL4K1rP
D84lT6PgFrEr7QCCVhskctAWROIcYtajm7BwugQP0LJDbh/3q924FYY2VJzIgk2kWPZ/2AW5TtHm
oC3HVp0jSyF1S7PfJjFValsAMMUij3Rf/2TeugUZRPeeriZwhyD3RBtGAeP6UipcPgoX5S0R7meY
2uUzOBP2BwXa2Pa+xI8LSkUvz5XNBT6X/drbp1ZZXfp5wPMZHqAcILQYeeQa58Q3bLFIHcM2ZZit
xnMOYcJx20athHzZBMxoFhbTAdLYoC3k9xfhnMG9YW4AfwdNC+5smPG9ZK7pUokqYoWIMFrNz/OV
3TaZKS1pirm21PP5fFfM0r4Ow0PGmKFGsY2wF7kAI90W4UYFg1SIBraRz2QeWz4K7BFvu707eLtS
dnAHUioD9UAYogHpPXpRT4i++8cWWMzHiCNtYa/7KAebGerxuPlYaIWhcqhv2Yfms5/TRAQa3Ze0
FKbwC8GBZs6CTcOAFDPtIsZzIRr0QjatYO8j5F/XoWG8LrzsJD1lLvke7lskHZB/zd1VJNUVSeZH
2CV/S/vZ9EIK1dU4P2/BKx3mD911jF6wPLhAapc9LbhTDmruPleZDdZMEgOBTrOnzs17/HvZiylg
fQr1vFBUp0dTbZv8shQ1kDdmyz5Vyvw0QaCr9L2HWZFxxmQJiVtLsRe55XChV+q3qc4lhtakJjEF
lBPQTboxNd88rWdLqJQzrVYZgk1BoZGtZ90OtdOip63JIMQhJR/wJfsku2aBzEUFtZEBKnZzxH4u
Q0YbtCJVYnqVUQL6uNwYjfnya5IhXCbF7GjIOyYuewSxQBb8Mekkn/gMC9er9jC0EhBHkxU35vy4
7qvZYolA77bxyhKTC4TiQG2SRCBNkviZVLOUqjg5n0MTQPUy2XNbQUaltX/OmXVd2CWL9sPY6C0d
2DQG/+IrOcu/aFulc8CVfGEaW6ERFCz71drxCKJoQtqR9LnAM9itUhv2VukLIdcBHPPuz877AUGh
mYIpHHCDHgcLyoZ0m9P3sePER7Gz0HstJStxD/Bq85oBNpv8tGH1GOa9n8obqo6CqJW+XjfXdVuV
YitO0yr9iLQtqas0ZnSNTOo6n4sL4ShD26upYzMxxGDcUslfsS8x6DIj3D0ePwIoEexCKAJS33Ic
dnZtbRrQPJFdIsLQEuFw4JKMG0W/hBhG0EAXWlfB2ic0491SEy2udtuShY2mwTV/xZ6rdt7WvCN6
aMMod71l2q7lZ8rLif8z9nk9UN7dTtCWOtNoBfof1WoxkvI4Q8JSEex29Jr9gQKuHNv7ospPd9fD
5jO8CYlNwQ6JRZxgFMpmaxE21ZvfOWWj8t30vLnvqvI+1zgZ9howzqbjYYM3Yb1z9PPFkYXMgRJv
Fn4iEfVF3k6++uqlb137aUBboCyAaHgHfQO11N6pfLrrgvQvmvi+WsJ0flE5uBNdi2WMawDRVSLf
baSH8p8hFYslkeIVswTfNSNsoyX60DY3Nz2J+ARIaXLs63QqFtKOdlxYUl3/WNdrNVHFlAn4WkRA
f3XjGbpNRzhvcnjPrZpbPrkX4uqT3ccNKvFEnVjdBI4eyisHz5vFDo+mcOhqI8oXRWNAGPAdFFBW
tAqG2e20pkHHr5f6xdREGmHZYsaJ7eFsa0XA26NsVWI+khsl0EVoVKBaiVN6IM9y4G+8VHYAnxfD
STNsutxrcMUcSvDWa6xC6eWciEHULJDUHFuuli+eGnRjP5C8EhA0uqxHXrjo7+Lyozx9zb8fsIX/
EazYwIW92At2PNvetjCg7tJcqHkmSTGteNdbC4EzHTLdEQyHObiCy5DYowZcz6c0eWDi5bNdsWEj
nsuWSg0yowRmNCG9HFonK5bRHmRxKmI24tbK9y0ximOEMuGUdThzjS71d4fkaZiQoSgPXe4aaQGy
jyp2sE/UjHBW8S0Q/78x71KThfIZDynY1Np/YicMKyjR0VEIntGxNsfoi69zgZYHw8Q1tNSsggcc
OgnglU+Jsh5miWPkNzI0DSZc0ELG9b2UsTsVyYmrPjggBVeRpctQu2lBvhMn+FkytAKIrR1G95YK
WATJk8qvO1k/4PbcuC/ADtGjbwpbnBvsTDNVrhe0iC/a9RQBgSdeqTPwYe8gxNRKDIhtBhx0RS8p
f5kh5DSWrFWFKpI1VXnzfvoux5VsXvq89Xwmu20xa391OzFeR+bXSCKCAthiJODxP7rzo2IwH4co
xJprfpU0t55QICGiXRDZ8ln/y3PHwvBFfCKUO7JWRhI4k2m6Y509+r/1M2rBp+Uw0GWI1ON6++de
owrMyyUCcAnFM5QMji9yzLiyvl9MMsggvF2NFOVTbDSpVbSHTumRgmywjFDRQSwfZfGaTYzvq1u+
0CzIs/CtRki+8HEl5O1GUXEC06IIqVBi4fVdo5ZiHlqPKd+89euCIxGg706cn0ifbdsckF2U+7Qq
m93TXpGeUqZ8ZQwuqW+sTYPrGlbYHW9r7P3NELNe11NPcvgjfi2p9slK/nZYVPK8T+X1do3dyBd0
16H5G3Hu07oggTug7QwP0HZFjQlUtaldhYdQv/L/+G5/pjNFvE4nIS7j3B8YLKew9MTDg6tJ6mEL
bNBGfigjSIwK2wowlr2yH8M3U5Y1pZE4GMsfwhvsKvIdq4tTERUDO9w7ctnsh5b9Thgh7QOJFUsw
qeboBbQ+qEvZYDfpLpXWGX6tPz0XpBNfn7TMSVJG73StD659oegU6gFE9a62rxMmavKI8pKI7Cjm
jr8E4iQ97pD35q1urHBTzqmapHwMxdJiphJIOReuX66jrv0HjPNtfVFONRr2H/M6F+GoprUoHEXm
dFbJdIEdlBYy3/K/NawF530cvBV4CmsJzK6LjW1WW2nflz3IhwtgYMf5tFfH3YycQeBc+GISq0Gb
8HY+UJ9nLqsYx2xjeskqmjGvqJRkFBQpJJm39MrAb2NKCPomkp8qoEwBxBvVGP2OUwOEmcGk5loR
YmyhqiTJMeFQd1b2K3sG7QhhBPjjmaMoxZ7NsQ1xWe0L4i2RfQ7+5cTr8UsRF/ASt/MfzJlmvdyl
iEG+Ho8gmcw066YDfyLWTbB85d3UaQP8b6djKCepymkgdDcl50V494cW8FwWnaRV/A+OY5yqykwE
uNFMi0m5vfVW4exHnkZaQ/G+WG9Ni6pphLxPnE5+Gca7CLz5KV2t8OxP+o4EpRk9BtYNCendXtbw
GeRoD5SK+jDHFmQ9lgEmqr85YefLC98YUIb20FNd4viroxtrrocFhWqvb4lLU5nDkQAkIY20XO88
K0iNPdt5zgZ5Xgukui7BbrTzJmbTWgoUbDDIO033jPJ27i5mK2QmXHrlVqw7XPYtCgWHUsyCo6tq
+Hc+vk80/fvO2KtclAEI5p4Yszb4CDRoHo6HC81HWcMNgRrh95jsjM7FrNaSoBp3OJjTTxlhBJz6
fzAcR94vbUYf/1qg+FOhrynvhU/69Zg/+QXOr7MmXR5Z4HjqiBr5h4sd0of/tvvjNu90Ui5CkdyI
n/SQ36Yyz5x9yfLocsATTatuUkZtPMqdPwjIMUkt5f0pz6HIF11Eg2fvRrTg1aa4zo2zKvARO/lH
QocT5u3ottlsSGsROZiQLq9q92pRfWXI/2dVIzPP00FkK2KdYRr06hIwLSM4VOulOsjA1RT0VJ4K
raxOaaJOLn4PIkbJsVZ+bnBQt7Y0cwebAjxqyZiAs92IfogQVL49U2e9nVTiKWYdPnmLHqQ8AC61
UNQgY5G/znCOsFWCYcIp4JYCTcvwFz6GjD0dpZ3YeewW+jbr6oB/cM3cSVAFJshXrFCMbDo94Y/f
du0gvbENTEiqNjlsDKkzABRTusfqCowcxiWOTPp/i8Wyo69p/GHzSKYy8G69mzTGA/ow6E8xmskO
uqHTHcp7u+4fLlEaouNF0rB4176pNZQI9jedBB/8jNrZa6eizVcFx2uETJwqoyzN6ajMdoUalLW5
AYyMEOh52J+FZxWeVSFq0DpVqvACvVRaJIv5WnU0nybOVHRVp1xTsU4iDS29y7bniL6iuw8WMANg
/p/EbsaBzECiIFnbQHby1PiR31cKamViwmVyXkR4m3jN5OL+DZbvOWmeCxa4/hPJ30HLYUc5ISnt
6W1rK2b3+BeUk2PGDSCGnFitrw6OFDmWiTfsWoUvyZA+fTTYLRiBJjXcmPOY/irkfsWV+Cds/r2K
pUh0JhMkiGxHUzV2FWuQNLWamQ8JBQrKk+BP4W8VE15lGGht+csQ3gzhX1LFO48COe7n2BIpGSpt
gW52HyEAP//AM+TH5Qtf0hHVvW+IOxCnz1VoFlShkr2Px7/sBYRUWgbLiRZjnxh3qhDWjPvB2bAv
W6K5M0dcgshRBPR610W+j6QfY42bLPE3M8yBJQgG05U9DgPmRwoUm4FXn5aEw0hOWZy/+MNu3mC0
dmlnLb6ivH+MUBO1FIsYiQeqrLtt5EkFyjgHE1rOAyugIGOW2EB79SNlG1jWvWxg3K/RM/UU2LYB
PDc/qsjW+0YO61co37kSAx88u8gvDull0R+HQhF516xn6HfYL8qZxO24FjPiTBRwfgHnmgscXzpK
z5YnDgJwpHC0wNz+AVacjuMIY3e92/7yj3mViZUtXDNZtkqemGP341JxCdSZnVArEvql0RlD2bnl
3WGmY9U8pisZIE+i8FSylRqELiVkpozTich134tlNPGsat/0DqxMY6ccoLsa9KfxVAzfPgIeZPu0
oGMBlPPO0HFRt9WW2N0Ui5oGmJgbexWSZvO0bY3+i00Anu+C700AnXjaZiLX9X+xy95ONplxmhL5
hv8qYUiztd9rfVQ6FydSoh03w3R2+qIYoDIQiF3cwFmLKiPREfj2olISVmogoTTG9v3ZlS0DPfJQ
Lx+1Lx1T0ePtIXjZD/5mFevfXNes94kclwL3GCL2bh505yxCMofWbaBPAh6lb42yRMKL3hSEIYTh
OTdlw0Z3+yFwTEHNya6ygQoW/A75CeJIdhhYmy9jcdkcM25OkMsNY/P5oXD/l08aRhSUUaHP2h0e
o9Wig2zEddtNg5Bbc44x7ab77JZXRCCKmjzlVJl3pwH9Af60UuvciR+nFW68UJ7tlU+3NSWwxgvd
HrWYlLuLqzJucTQwI1jtED9RvstgUQ8wTeGDzTMLUTYesxX22DFcaQ4BUMpCb3oC6ogTU4TidRDr
XYyEalV8lpQ7t07dVztbr5GQ3NEJkGmWRCyO1GDKTq+dSBIOI2pMKLc1fig20SDAd+4JB7J4Od71
AFucjrWzKH1sQBRA8O0ugdKFjpWyZr959GeQWMqZdrZmFMYVIKOaCg6vSoSQNy2liWr9VvBpHztk
nq10G51DaGX30nFTsKg69ca3nYJSzyIJdaATwbhpyfOf8SzDRw3AvyCSSE1qWlCStdH8vTFzzjt7
CafDfodHjxUkzObF5oKD2ufcnyqW2vQo3pwX0umV62WpmI70Zfj56w0j55t30YSdm9kx25JSDIC3
TqtqAyVVvF21EZdXl4CzisYBVpe0qpfQXM/WO7mgJFyq/F8oTRXvl9Bh01ILW5scWtSJmXzFKKYr
2f95bB36ObMEncwLR0OeL7d6XV2QvNXibEAcln10B/CKicx1lQwl6tAkGTSr4GGAwU0+ZVnzyUFR
DuovHzUuxfijUDDLo9YENsjTnUrz4WYKgz1E8cbFecDqtTJEK45Kj5LTvB2ZzKGqUz/IkX8/aMK1
NGkJopNv1aROmQm7zVq0zVf1Ma/XcpqBr/KjePSTOl0KFH0Z1xWwbCwX1JAOTkamE9gUnq+qlvdL
4RS7rvyop6/qH58J/4l5LvZ2qVbqgJEkHsY21obGqXEWep2shA7rQhQ6XNpuFrPDgVkV7JUjnutu
WvuXBQcdZ3EVhqMZRi5eBtefVH3SOqVTquY9Xl2t2YgPkTr7oKkYbwxQsXUNrUTPfyuYvr4bYwa6
6FST8BBKQAowqCzLN6Vn9GKiPjLxa9+icjNyT1VbEnqD0CO99cqXrLVjOnTB1KpffIgIwvHovcNV
Bhl3XCjCK/InbTt9VNP5Sjcj3lFW548+UXFTMDy1H04AZxiG1tRIjFRpdK614mSgElsQc4Psy2Ck
yQNRGTeEcoynMEiCSHpqxmMkc59Z5c7hXRTsqy/rRHJuuYEHi/aplB1+LiV0ar8ODOL2t2V9tISF
4S8SPwxeKftaex8Sw3Psl3Oxo9aC5KEC6iBitvjrI0d+G6Olu2VXCdXINzEm3bXkLzb5Zl9yY6I3
qFgNx5JmoVsBQ9iM6gRQd53L4b6dYQQhoOgXS5ZlxQFktUT3VTpR7Z+GZ4EF+MjWeZ886Tt4lpcM
XcyP9lFY+hAv6b5YoGOpHifNGJ9ZJisO56X+EjDTS1LaH7JcUWf/50J2voDmHGEtCNkiRYDYIHw+
mA1cH0+J6k3+tnQlR4erpF8rb+VWDpy5x8umScYs0iyhz4i0S1wZQ8bgPAuz2XpvajBEAQuF+4Ex
UOeCMMXD3iAF65XTqN+qygNSDDEd9kmGUDtPQPGcc8SSPw3pJGo9sob0OvU9/iYXHJmhWs9tIhW9
3MbR6rdfdbiwnM3bX1aJMSyQqyvghIsfSMneKU3j7vyZB+6xgGyveZWayEH3qWWVNIVALhvsFXb4
M5zN2var9rTrwByU+2A6TCymBATLc4gLH7u3gaWPHKaWXkQ4GePr74KKaW+70SSLuel7bVdkS6nk
SvSsXcm+b/UALCuXNZsEvYQn7HDkF4yHNH4Ewt0UVIEl6ixROXk0tW/XWGH+vOUk2ePjkW3qeoNH
cxy5T1n1XjYxHhopqhL/TcybtN7dNSeYWvG7aDYLgg8l2BwrrxH1GTFZcGyMgJ7+TK9x+cZAnuR4
pnp4WihlLhFJUt4GSVj/okzjyk5vDJL5qMJfZv9yp0EFxfVI+xYwNxe+dxCN7Nan7PnnGX1jdThO
7tSwN/MNeWGRdUUBfH6Gmk35GOIOeIY4DqPMEt/PbbOvy1CztDgx9yHI3dZVhj7YXZGPi+O4lJ/6
tHGcj97UBldVOlCNgwPIq/2+MVu6BMXFMd6pxzMj0/CSC5OoBAtLkDgu5nxcrB5KzXmynqLf+XqB
OQhuw1ZvflbPXyBCzJ0be/XPcYYyDp+T34MvYRkK+uXv2mQ5FjGARvoc+ol02FbI52+U1EApONj/
am/t36T6oEVAG5DoHOXr+jfAK2GVwwk86zlDq9i63US/waWxFOUgvYwI/XXuxLa9vYDUfe7E3imr
zY/aT8H2i3T3RjNc0nCYY619cWXlyvqJGzuE1dDKRPkkfvUG9lgimGAlOdqvFjTb+y8rlCN+BpUP
eX4DsKIRKcDLVod6xhpPMjkaJkXcnGS505MEbIqkk0u6FgJzwxvIWjHKFF5UtF8ARe8Np5r64mGc
JeBT6Qq7+t9JOzgHOI/oQZfJBEUuj2qZcp9LcBNhK44VhNwOJXLaFNwPnLaj6Ov+fhF+X/t+rsUA
cyoUxyiZjuceR+4Hh3GUNrL7bNgzllSDaPK6JoHQnKJoGC3qBKi5McADLi7vlWcETdvN/clIZaSQ
8FK8I1GlkGw3UhacXGhSsOMKpVW4HK7/nO7BnBr9rw//XCLrpcvnbSo/iFA1Cmm7400D+/FD76Lb
/nn4vv1ZxKRPq8ReyxJj1bS2ZJb2POQepEEcCsc96i5n9wz+3jhnkibLWyOsgRPsMQgmr7ZRnGs+
ljVP5oskMebRcmforEtqnFAl/4vv7tvlVfhEa8wuQ3WhnScKRSb4ud87benNJr4puQbCv2Gy5umC
lACcU1RkkyDUGWWlsiKAdXlAspniKQPZyzZyH2v6RQz6eVdtWgh9pUOAyhynmzWLahVUHHNCRiJm
xIw0tSZnuZRIfRXWtW2IZc1vs7hg/r1ya8zBi3cQcSjKmd+ouo1/Yen3eda2kQ+HcwLLU7KMv5Z3
3dO9s0o1wj+GbCcH3JPEq0rac/674ehc2SDUEPKeuISoF22DhFYD35MemuI+hX960Fm7YGIVtlEL
a9I5zfjKXIL8xSe76minUWvJpyUxPEAVUY8EHPqNRDvePOo5GKydc3Q0LmSkJnWGElpAbJFZFbwh
HsUl/bUGUBpQLMZsUOV7F3CYTbFsjOuFT0hLvshLXu1me4Jq1KB0QFkh++LUlz1fIdR79LveWurv
8afiLvSw/SeSmfNa8a3WoJwgl5rjsEr0VPjBueIxZe+3X3wxC4w+oR9bj42qxWFgtmV+7fyZBlAZ
+A+GPEZDagJPLl0OTP1kxEUWWjkU+TdQRmphd5TAcgXqlztN0NwemuHYHELQP82mOxhDIU/vePsk
voHIPV0NRvAtH7lThYY3fiXtSsrpfEIaTefnYOgD0ELF/9Lf990v214dvrWj7R5UZX6bXDddT+Fr
hGzJGdbthPLgOz+gF7rmrkMnu/zfoSn5FwWNytepNrih4oOZDEgH90g5joEzxqYrwpC8j6aK9L0P
oO2mMTuR4VZs0dKBoi8lJbgM/p+byCevVvDLb0fHQ+rF4v9BuZaBEa8jENK5wz7bSjr5gWwEorED
nKEToXFKiEYTLlSjkHhvjoT7l6mbWKUHGSQ/HVp3Q0kXUly86VLjLziCdQf0wnqR0n/7M0oSyeNO
IE5AF+s+hqFQ9754G7Oic70mRDAXO4b4Gkyo/ZuWcSHsjj1Uj6jEBxHXGsyCJ32qCIt1gmIm7nWp
dsCft3yUQZrK/qik/FHw/n0z5IwZM4NFfGdnfRybeQI44Pzvwz+gQjDQ0LsxD62wM29L6IGqYhXM
n4vZHtKros7JN9g1oZNe3/2sl82WU4sm15qUk3MMwXhgRFa7xXUdhF3RsNhNBjFlC09rAbrO1YU+
ve+NO4iFX7EdDeJqc5LonGgFelgBRTPtlKhyUDHAOlZ6KBKwLNsAo1KU+H89g+BT73gZ7bV3Aooy
d5JRiKkY2YntUQ6G1k6wWYl8TpZ1RjN+br5VhT+s6iUKoF0Q2WmPTxkHZN+g8NUUwQDXLoKjhOp/
o1k8YfeonEw34o0LA/ilOHThjoaVG+pXroD5Sid0rHr1lhC1y6x7ozxCUt2vxT4mkFmk6uFdwpsB
EeYICmrKadXI/nGSyXeWu20uumQ8UELZc0PJ0MH9FKxQc45C0F4X3DGx3/KAi5FB2GJ8snt4uWiT
Z0CWCPzWj733WGt/P8jvBdmr2HfIEfix0GhP75VoA5GVxBTKuGkuFZ+COr5rMzyijrdiiyRYv0LM
GmKJW+iJEZ0JCl6p4VGpsm+3n1S2Y6r36H+Zz6JFjvMYBQj00z3UsavBTKeUn6rMIWgEeLdyssVa
921Keqz66LDkNP6+aZJ01N1awXgxRIzcleWVne14vwGF9ZcyXpkb8Wt/SS3HYLZTaIZYWLswDHOF
yD1h/hR4wVJS0hq9VxIxOGdOUUglWjcG/DAfhMILU/grUpwNulmLOF/gj3YNd0J6Ax5+Ga/prJOH
bXA6Ix4Ne1hqSYKCOt3oZNLIMjkbihZTFWICymVPdlnGQmganfZhsWTJYVc3pq+lm4s8/Gn6/9BV
fAMuvI+0ImIzQnpuCd/Ckz83OngGzN6hT4skTBux7Eii5rGBxZMoeVw5WhHTKPJNk5h5M83ZTuKZ
zPC6QqPbxwLe+zJrYNro4tD0wwGEpgs7+z8ELbJ0tmpGcTKuS0OUx429UQ3hnybcaiMIyv3XTiaN
seSvJsyXV7CeCzp7fHBcn/O9t1BbchtU46vQEyjYHWmfFXEoAG9ODK8MbcrexfiQQbPVQ4fm4KCq
5BT137E0xtx28VgoAP4nXRg3YyFxFGAsz0EMw4IuCV+0tLIkOE3pyr4kf08HLSQTDwbkpvrywDhM
VmNwFpB6xh5quqfHm1HjxhBBX00mUVO9JT28uE16Dgyu0DTccTqkLC4DTRyYj6Wq3rhE/If9Nww7
MQdXIvhqGLxyNrtvAh2+8kCFAalyQM/KV8A+HDenmf3d+q6ZjZY6CXUWZyAT81Ft+pHUXb583rER
Oh/SMlzpLJVAmqNBe+vL4unjj7GUz84YTAxR7DHIoH9BGQb3ys/CEzLg3ta34u6phI+F2VpEsJ6S
+DGHaDoaolf3SN+WR7cKc/7yyOGqwLmaqe2TrHHr5CKzSDijhL2EMrJCAZ/dAxRxlEmFgAtI1uwc
bI8SeA/cQgHbcxmPCPHuXLWmoTpzQvi6oVzA05roV18XttYnlUG2A4lKkh1eoyP/a4skwGakEPiO
XC1vwpc25zL3meIeXsWhB/RM68cor0QVtVZQBW5UikDxmqCfDLUSftUpwkq0dHRg6f8SSIEAjf9s
4lHR6YfzkHVQUoYG0mrD7yRBQ9ao5sgKTp26jeJjHhQNz12vC8bc0lnYKhrF0gZZsWoxdN/L0SO7
mcGewmkZsSlTjlT6zkIkAbX+saZxm0dR6/EwEAFSfB6Q9ksWdcpHSVdDAiodo4dWp+SoJpwhRC4/
687sX8+Q8KAPQHUN6VsbBAoy70SRq+5j0CjnMLfiUAGjHs5A3MsExba5vSSj3KwnlMTsV4510J0h
Gd8jSkuhL9bvBqzHYcmVnGWZ4dbYFRDwfLKu6OblcYddN6M4h0hagXnPI5C5D2DRrBVUb9otaVJb
/vkUy6BTvHELf+Jh8hjnFFfew5G++UDLNCqA//ipIGILs0xQBHqQ0RY/zFfhN85ko2EHfb9DIJZL
pl9eIZl+z7QQO2mHi1xptAg05rwSzKDtHUCn8vnctXsZo0NVSzZgfd+9RIhTvEKJxynmsdM5QV/9
zFO0sWRNZv84kcZtXJeBzXHdfdJMEiWllDr9FPpFqSTWCdjGyzSLdvXm/qBKD3gHTxaTpuNNklmx
MOqyLSAAGj/Roz6gX1wCaM0Rf1Sx4ujk8lrfcAJIgEqD/6s59YYlihgQ8tTViMZkGUpM2LEmyzoC
udfwCOjLGXsDGDw3vMRxsv5XgKPKv8b/791BTJ3ZtCZwS7F+A+qKe67nlslKBmq1u6T0r3UP3x03
rwqyPsjXYyyeX1/5MnwW2lgcIMiimQjfJQGJRj+0TGp+FQ/qts4QH1gFIYixBirKO1dlZ7qVNHXc
S5O0XKiAE0XYXPFG7PpQ2EVRTLgjdehoQ+LDrzwkEqJA8L61N194DY6mvYRcPvmCCclMaBORw3dt
1McyD/jZYFkdirXPulb1wXJW12VyuoomgWJ7VuNuyZxhrkD99S3hB+6wqH6Gi6Yazk4T4uKhucHD
iEL93cag0Az2Vv/qAmnD/mCjEZeDXfQEo/Zu9ArhfdhouEyfPpYnhJhwXbGr4A40OHQ9FH6jr8Ti
kenaphwUuyp7Bc1HCzFVd3QEoaTbXqur2CM6AvWGagWYM7g0iNQ2UsvjEtAUK4lGyoveIZo0BZYy
HXfDN0qEHNuAHmsa0wkMAnIwsQPRb9BPo+YXj4LAE+2QhCtDvFCWOWLpbK9jSMAsCBJ3agpfAdvM
77aCbdw40tAVGP2w6LaI0+7SNz0mWKOFhQUSSHY17v1a0Odsj1RBPq6canaLFyXK56raALYD6IWT
X+ULEhbBeAXJfH6lnWp5mZkqzrqnYbeWn1UBT7LApucLya7v+6WCoqWclKpjtOANPXpMCtCKzRsi
G6mscIdVeF2AgGB9OqI4r95d2xMXoreWt6s4ks5aIWFLvmk7BONj/qmklvYVt1LYiDx/HMEu/3Ef
9xTYPRo8McZsZkzmqzSbJlgF0dYMvCT/er/sx3Kpt3z6Y0jLUnhTG8sdMy5U+OkMcme0+itn3ISg
lciwCJ6Y7PZyqN8TcPLF+DdFD/kVWi/zqOGwJo0iLZbHPWfjUgFj70zDiEHmpQzBTErV064qyboA
RrRpl0Qlzjy8actiEHiXSOU278v7uwgLnzjiv9J97Uj54jLO8L+wrq9wWkUWkUK0wkafps4EsZx1
9ia4l73TYqvLgTpCAcIMfwccu8DKFOrC2SKRbrjylt0zeHtyoDe2vWdMlIldkzNIq/1TN2s8YF9/
ETNdUE0/XuUWpKOfvJvB+syPpA2ut9+IgeSYIlC3v4hzQ9wVmcn64Z6ZOE2A65MFvGQRNsX5S7hU
Nv4mxtS+0eMwlavcan+xg6U2Ye7SZGUmBH0zStq2kXvMoC0SjOqzcpyVQW7PuE7TokAnbz5H61Cr
rdg/RrwxwEfB4+l/WXnW45xphIJEwP0hVK6euNYtTfFV8R+fekmkg3xmYXbIzM9zv8RdI6Ww7Ptc
1akcgMNqApqA6nUolx8XAGUNen8VZwkDnGsF6o3mRuPe/4RyP6swT9AgGWOMhIwJ3u59xvte9C10
sDkq0L+3Gqhv6/VmvPQluokUiaassbfD61YazhPImE5tD7zICqKmiImklS9/nq/qElJtmxK17FaS
G4Spp7MIvjBU6ySGwJgahM2KGUCCl7cCS4NT/JG1Wp4Vis8T0d+BIfeHXPyWXMyHqqBQX7rdeMC4
VMVq5rizAUQb8iaw6TlLmkYkPI1ISbw/icw490hKSS4GNG23gWBjW05yaqcb/wVay/6QvpZWutfd
aF6aNymYmKPoPlM0pdJMz9PvcvfTwzjXbs+MNm8W4feeJbJQTIHixp3xXD/WvKqoIn5lv9qhL8Ty
Zt8MSRp4esqtFfjbRvnPX/oG7i/4Jn2k1SLH9c0DS/dm5Cg2/FEyhUueFhfUUBbFQWY0uWyG3+10
Tzr17VvDRxmocNzGnmKQVSDkAxe07c7lJi57HKJHUpze6dd2z8DiDT4oW0QuFivuvQ+y5bHTKkoO
jWY9Viu9a+bybMATxLBm5cm2RRDSv1ge6FWg95NDS0oGGEVo2tLAnw65YVCJGA/th0FKkwgsTyqZ
4GGusap6hkuDEOUIsFtUf0nvgeZ0At85v7Smq/K2ptkiXc/Tf+EPicAtqVgF6qm9QGcBKaRPA3Am
H2TR1u8GXb0U0EvrvDXaJXs9k5TKK+kjk4U6+OPu3ncBW08MLTrHKDx3+V46UnYSPHQOubgJ2XBy
fjTUxMMivNJ/lhIX96NqiuXPNNUwl0XSapPjMUqtZR0F+74CWA1e2Q4dANFc5Rl/jrWFdpV/gk5w
ONCZTd+2gyv71GVwvrOp77amuy54XpQ6QCWkKdZIILqc7DEF1Y42x1evGmiwWCtdIkt4f+Ac0fOQ
JD7oS6gnL369HI3krYSeEzn1jh4N5rNk9iTIw7WXZc5xUJkBKI4U7T9NbWxUPV5USc6d9Zf8FiP5
WNA74a4g9bW2LNGhOwIeuHH4BWigmz6tIIDm4aHyz+ElTMNEa/W+WDqj5GJTY6ko61piRRx+5C6S
z/khi7fKRsHmSJqfugnI5ot/RmXRULGd99Qo+XBrE6MLnxhCiFMCto3eO7kPiE0TX04aCakJRSXr
XEm2lB2ACsNxUMxxMTsxoPeM6ktqmFcaBt3wbioFP044ccudiWecxPA2lmWr+4KM4jHntUDb4eXZ
GMaSEfTB7olykovVD2AuYeXGT/2spa5Ni3A1IV38+pW8zghRKHn7tgVV1Jx88vozwWg0ClOyAzwk
fEc4IoifTSZ42pvkndDqUmDbPthaZ5pNl6T2oQolnABoSSJsJv/vOQzoQ6lDrA/AxJvieKjtHVG3
oVXyAPpWGggcoBf0Lg5Q0NoY7SARAhLJLouq3zxFC44YaCCMGbNq5XpAS5jdMDipZWEI3UHijjni
Qqq7dvSzRKbuN18V6dtHKlbhAGxhBIzGxy4D+RubzHg7Eu8Aqf/fS/3wv0ES10MIhbf9UgslW74Q
Q+ieu8bIhau9Ua/xxEyAyU44l6ErZde/N+YBug6NyEP5RvcEGORvMxP+cRU9YfD+bHlflWC7KDBp
uRkedfWWeRlqxKRQ+fyEwVzsTIVB9sEOyGOw4RCvyUfSmZJXs7nA14F9hZGCTfteZ5dFT7ScuHXf
Rxj2Xe6mHlAtlxAAAgpU1l56OPFECChRBiIIIsytJ4XAOt9LsB4h9b3x7KlV9V7EXnXSQ4h5DCXP
jrQA4/OT3I3xCQ+bX80lK0l6L94IgAen8ZmtvSx0sstb4sXy1v2/PVJRmn6dzzPxBukHHoqPeyoK
Pv0yQykr/S7GiZmotzjY1zLFTgMjRdFvovGZcHOFNBTW2LNWB/x1EI+MMqg7jQJEexKExdog+/MS
0xuMxg/HxpIX+4/0Ocye0T6I1hUd4IjUgeuDOh1Px7SYIfsdALkEA9Wo6UhbMATbFKExqWDDCvIr
rV4LTYpapZgb+FNcpPIjeT+mAAH/dVuEDIHVV1LfHXmLyBKsGZMN3TP5bZnN7kMotAw0wb5gn1Bs
RYe7iYyGwR92aI9AE38/bEX0nAlDBOcYV5Rl1Z6ZCIHOEECD0koMDNCkdMDUsJu4Z7/QH/R0GQeI
JLoo/crK6y2knfgJUrWk+IGW+42LFCc7MP8ejYa66MOZdo9qXhi5jrziBAlxAlI9kdHXMJDTtIO/
bzrezily/ehmTwDPYItLZoZ5XUgCTwHGg4c54iBky5/1dtPBKtGMANwtK53PYjSC+uUcVk2G6NYq
6AF+I7nlImJvMi+RNo+CemxuTXP7LnOpD92MkKNQAwPm5/mjMRa1vnGytrX63tZE39wXw9vBxw6/
DLu7T+XXm/7PjuXqlpKgpTS951eKMbo09D6Nn/dr1DQ/TVgN+8+fwv0VtV2HDZrvskU1Us3I5qXD
aVhFMDpv0S/Q8WroRIDOJ542AD2Ol719ckOn+sYwz26JznKlVFsUdnDGiMWuzm9hFds4OtA3UK/q
Dl6Se8htmmWTdX6vVIGsmEiGi7OsfaodtzvyLEhuE5ynpqZ1rcxweEpwhFwC3AvMuP49Xpi98ptr
+ggG1w3VGJSasQnkomD8M7EgkybSVXUcepaDi9MBZik+8p83/hqBIQZqQYTjCvS/4CGt6cdPZzII
vQk1Ex2uyipfG79kYTHReIYerMDZPTOtrsqZ9W7gQ8ZMr1x6bHznmDsA3CY1KoWiY4KThLK6JYds
s4Sg2pyo07IXcq54j6jme50f/QlLk/z50Cdwc9McKGNgtzlyl3RZyha7UW2mlbfwrOeKFCBbCxJE
dUqbQw+suMNk0vNay/Th+zwW23fjd9M6S+7xscQoEUEZ+uCde3YNmGlEx4yDx8C9Si2xJgc6qHcU
ILfABZEetYzDlXkRdypgE5JSwh8CzxU+ZSrSOae5FFlwoVqk6jE3vd2VeKlUHKFAMXO1IJ+vb2lR
pD575Uwbs7ajnAF0qHlkY/ztIKhoM3+a5A3AFKG7Sqmk8TDYG4BnuohmcYWOqyT0Kt+568XhmUIi
2wqou3aLYyNZAZxSUazqnGQNvsmxjPQHPERpbVOwp6VNQOmyrZXNRQXmhEQ3QUJWSS1G9Sn4YZk8
ALNYErGaP4/hOt27xpRap3Kl28uYFhxWWcX3KKzJFONzd6EAQc9NwP1saY6rbyh3457DU9poiwLo
gGlMw/wvrBugDRuXybyfcxFfKetjZdIL0Mszk3j12Yfn8H4BVMqvx48C6kUv4RkNwwFtzCOhNSiK
kd6rmWiQR8q8Ra/nyuq6uZjfeJK+uNmQkLfs10zEbCRg5GXU2qwCkwoQhSw6r08Zw8G256htIJL0
uUyDCIGym3PlgVG1ISPuKcZzMGyjTYixfKb0TcXb3aqhOvUNUvFwkizuYPeFCQ0oaN+PyOTyUKms
vWljTYosrjUxUq/aUXG19hJUEvIpJ1lAMPVLSl5NYgz/jXZvWcuwn5eNUg7pLLW2ZchmmwcRC5/K
VQiNfzLppQap7Jpnwja8GT1thRwAdOt6+tlcDoEfV/WvhhJbqEsPKW8otNVawXZeHCrv/7IBxBVs
kUXgDdYVRFom3Xk+6HUIe4MqviOSx41hbrBtc/IcE4U2arDxxnVM1csK8baAlvSYeSHWL4Ev+E1U
RZC05sN23KFSDpbWxZhb5wuzM3Zj8cBpE6twOO1swnC72Ir0/fDWMqe7oymqzw20z6RNYtbjMwGq
6GGOn1fdjjhT6fbFDjeNMXwIYzE1DW47Nhd85fao4BqOZx7RAtHP9vwARdERqRn3NuPMIjzIDG9V
wcop9FxLgIVRIcE05x9p+PwaqRHcpvnJcYzlrn348qkCw8Jb1ONFa3znXYMcIvZ+zMaTXJws+Pq1
VgDe9Mvo8WtCvFto9K8SS/rGiDHljAPzvlRrKnvjXsj2I5vrzBM5EELWvTuiRjVdMDYayEDh4k+R
E5XHegCTcmZw93J/QCalXBKN21FmXpD0+FW+me/0KyHUELTgOANP57upi44OmS/rnsGGEc4Fz/vh
IBf7KCzqMd0iQ2IGoag/YB8bRGaLBFOcy/gCmKOjDPPUTBBLqt+qR+p0milA1BHitEb7vqPIx1XA
L0eyywMCNQ6t3HqokjYj1gxStenekvcP13UEZWrR10vUqRFDpmPR874vEn/ndIWHncqLDrV0KUvD
l3nd5AhuAlAsKCBN0PMR+k9Z5Z8cFgj98SKHL8T1dlXSSUvN0OFfK3juqbN72hVT5Xj5DfKEvgXP
1L/+C91wEdPTmxlUaTHLI2vx1LWDsi7rSk1XnvT3A84KqdoD+r+ix7x5jno/WfI9sFzc+1bTWUvc
/PU/Daznuoy1kf9lO8jmtQouEPszQ5Nb0FpL4ddzb3ckEFbJP1A5lqKuObJMS1kmewR/f1VQb34e
E5E7pFrIVii8eLzHAlbKKWO+jRBWHD9kt9ESUxRlbhgnMxPxGUjYLHZECgd5oPc/HElU0HcDqP/P
62+pdaroqJnqYgcdS07cTOlQA1bxGwfhhfLos6b++bgRcEdjHhGw001Wo0kZUnIoxAx9Jz8sCxLm
Bg4uMQuAyMXOf+p7v2hcA35YKJw4AHK9RwxrTpOiJiayxTYA8cYVWhimAyPa+mWUH4SNOh8OXckm
ira5DMj3oigI2H/u7z3ct/Gw5/ktE4eZ256BHj0V9gICnARxL1D0J1Q+bCWadoaAaLEn8AYMXDqD
0rD69xGtPzkYIvj9NV9p8PdfgIkEIn3JxLzet+WUQUJ/qMnjtEOb0cEwSvBB4eH6t9m4jiuu6qWI
9lYZJGumWHJEGCw3ejKdrpCa2CTkBy+PnOuw2x0WOR4ibFcJtl4eYj54Ik2EYt2BpM/b966/agnU
HznPXiVL0FtP+VMd5Fw2SjkyiP4VOL2lOSx9GRTujBKnqUUwWdl3AEF+atFuY8vg5sO0zQhssRRe
EvcJrCH3jI5Lvgykd8EC8ty5B4g8uHeli2UiPWDoKs1X0UQK9kVudB9TblAU0U1kUNOmYtmFc/CL
IJXkK4x7/b2QkR06c96VESlG2rhppH6pNx+i7vaOvghxvIJVaED0nb2ts2gx85sX7u82oC6CLuzz
PlxBsVEiu1ZHC9oE5CTFHC2zYcUg4tagnSahJdUhEmcgRbIc9RUsKzQII+UF9RFM+b8jCULNn/aq
/bLHXg5JiXjnG7cXIHAzNKxrLadqoqdMSnDv3GfTW/RwubcfaLPRbkAvKkRbtI+Wq6a+TDMDv/G7
vlt9iwnIgLTeM2hLqCf/cfUoB0+/FKQBJHPbk2xXBD8slTJi1y3CEPFjX0f1w1U5eviV0iwHYswk
KnJgmBGHj2m58TDJl/DsX3Kasi525X2Ntlv8V1dLyNBJ2VdPBSNRP0E120VxkjGepTeE/WHV6xyE
9f1SOWBC6j9Z6Js0bhhwVkafEv6B59l0gy4LdpPmd61NK7I5oUvD6AApbgrfu5rCd0V422VorGB0
62R+0B06e5732TkRgCgjfFNgp9KVyMa/6lF37SgHQIheG3wU0iL2oosi8OR464ZUjMSb2mYIHDDR
Wwy4azZ/tHetVz20XimkMxmff/kxJvcjkCda1jO1GxacAvRB4rFl6UN1shTvHAMLXvf4yCLOTMVb
X7BQqSYcFGGebUM9zxBCMJ9LfBa4NVlVVBKmQbL0goL4hoKe5MwwJsEV5QY3AVOR7XeylU+m2hWj
I+gPkvHVH5fwbsiHArjRM2vUFlvyl7fvVjQD72kp45Cv7rJPyUFwxeaLa6MGXHre7G2uEcHatyNN
u8vtqbg+dnS8IS5NNTrwQMLL2KSb/JL+vJr8i9FTwAhF4H9BfVULMtsIPVU9KGFi6CPeYiQjAsqA
l2KswvXTHfXgeixsnIke5A96Wg68V3kLrWaVwv/xXGh7oY3KAyFlbMSM+8DkXj80xY+Lvl3+GyiT
Fi0C8x6C8uENDD8SP4ZWqsUxfr6qSaOTWnC93hdn/tAKVBwvVyR/OYC+jKguoeGZQogL5fqXHNmb
jK+9LwUP7psOotHJtDyJbKIoa3t6WaT2lESATX1UZXw+0EnWG/uc2ZFX5pHJaYti36405HYV01q/
oKUW1zv0yhOxSaF1JqtPhzrn39aPPDluVawphXKSgByT/+Na+/ZmZNrFGbxaR7/JX2HP11iwFhMr
7xKOefTOjSQql48d2XhxggB7WLQMiroRPl6Ogbo31GKavCAnaIOXpsic+3MysBEnptCEJiu1nS4K
P5CdQkqnCYUtU5CfxvnRAJndbjIGSqaV6hyF5spP0F/KxYDhDm2OIII+k56b0T9MIfNxqxfSU3Qv
gpdBGRE60tTZFZ/11W82FBLmE1BBS7fQl31R7q07hgIIzcjfesPZtSI/HmYHdlGuF/kgtX6hQors
YvGv0G1j4ORJTGTCPeCSMlC9ovnx7IU/oKw2kZkY4KwoFMvzeuwcE4YZCGaQaQvuxs3JGVmuT9uc
ugk87TSE4Ty19r1r7A50+0hH/K4zQJut2ebn0yJzXQ6raTQpV8bYQliw6TsqFMhjuRlUSPCU+9a7
V26ztXpIHh8am/Uc+U7WjNN/JjtPOibDxuR2gDUeBeWvWPjhXaG+gB0wz5TKCJDN/iZXNYLwoIvb
owPR1cl7TPAz8URLbB/Q/Jscpm8USsVkkjwQ/tt+kG77+PaVXnLf+5Ta2oTw4NDAJWrRFL1Xu3az
RQwy0KU8wpycFOa/wrEsgItyh+ufsnU4cfFq3vOWWp5TTQqBcDfMoFEzmC1yxOway1Ur4uP8Z9Pg
z1HjSZtfhlBSPaTlbZatXjUtRD+00Q706M5wPF9kTYN68/jADyFhbeGeEP8C9SeP6zQY1NZ5c4A1
NTXGrSRugQBn2chlWqWIVoXAnjIeWis9wBnCr7i8EraDcVMlVdgGFrgTwFa2ZdEnONe1i6YqQrGN
tQ82ecnv1X2M12owCUfJzqWlPG+Wx//JRbOQFrjHs3jxOucAJwtgoTcsk+rLPIxRdhIO75bCAbpU
9Ez1nFQLU3EeoZc/o/3yqyF8ho0meOYjsLDURZAC9y5tCaXGsLafSF3CgIKZgyrYavUVv7S4hgji
mTIDRoHK0h09fMptiLHq/ZrYbq6529QtXblSqWqVGsyaKOINerjGlgnA8FhPhAzCFd07kim+Td8G
xeMjnoGA9jV9CTix5ZlHsULZcCYJWvTD5uEx8kHreMQa+UvnkMSped9VdtZGeNKDqr3FWOUledxp
oMNaeWDsiJjZjnTNzZklHvuIacFTeEHqgXAO3ML4tzO7K+7cX52oSXoYDMmQN+YeMnR6tdgaCuWe
JGSzpPcHZGaeeZaylgZ89Q1/eNtPbMxh0jv771UUlLxsUPiyF9Dle3tiT8YzMWR3SAEv1Stn6Du/
1/c8VIggl1iXYiMvQBNWrlEJqS97qr6yibuhAvR49sPOCVMWQAnO/0c2gdvXBZorYSiSMHP5DJAN
Yxg9NRgPnUuXZ14qFnjZAv5ZZQ62JsFnEmK6CSqBpSmENx3gLfJ3PLqJjXUTWEB3FjsPdoz6ikss
xecTbbh9a1wqfOPzyHrOXUwbI7SFIYhR7l8r1vfV1LIujmVsfzHHX6bVRa5T8yCJnQCF2Z7HtJB1
tWWo6H6Euj5brLRNqLaunySd7Pha9Dj6Y/lbiDQyXQDNHXi1v9UIBCElPzNo+RCXFdzKv8gfRpsv
VnxLw/Vc4sbrQWejYR9eIH4D6/DUu7BvYX4hYS1pnUZoAu0p0kJ1J2L46N4AA4lKNPoZZWiKp+oS
AwblnsK5EEAVpmr0AMI1m9b+FvjZnpYBKgQP0TQmtSo7q3hevkGcmdcbyqilVJ2rE2nZ9Boh+714
I00iWWetgQzwT7OLVWeLae/sNJ1l58tcwahCtnBpiuL7IWO7x1A3AdiWyIUNiQ+2snLxMh3QhdTV
lAcbm2u2NJ9S9Y98cJCOBc872xoUYZhVIA+1hke7KupNGBxQCxOsG63NCJroTYaw1O/cgZyDoPhT
ZGYgSpAlUI0f2HkYgZhBW/xGzloOksFT0Hc1sIk9/6ONxc3tJqILuYtairXmsC7A+ogIyxarsVp4
QCRrxZakhyXGQzf3/O/LVWysIiRGq/KrfUMQs57FBgygQIs0OPdLPh9KhJz7BSGruBXsevbJNnB9
ogUM/lZFYBJZcnozEdNX12LgEEMjdwXRrYfa0UmPWSgs4Qf7sNxywsXxPY3Q+LPNnSxNXikxk5kW
o7794rtR9IDb3+CYCuy4l0fK4nvkJhXf1xdGOD8lbEV9qQmp4eFEKGQQG0H1IeLmarfxb1I4Va1C
npl0ZzWedq1qcK2Drp+SI0/mf+7t/ckSnP+Ug3vKIMLOT/QoO70bpbNWmWDAUmhEm2t6T6KYt3Hd
oxQl9fOKx4WHLbBlH7eYLbOr6AJgZQq0mSLKzk4CPEw4bNcO9U1FZqAZn/gIaF4NA9mYsligziPJ
B8ozwTddTrBzgyaQvGD+aWWoYhqgtIAIB8ax40NaZoCyiao/K1E9gLD8Qq6WpPBQqFWLe/jmyqZf
+g4BYxvKfgL+zNITAwcm2nJGReYlKU4FG7skBaYfIBLvSOHEKBv5mqdRLArX7N38mCciWiC/ukpP
7EqTiS1mqoC5aDIU33PgUVoYITcgUUBOZaERf0t/D2xaJj97xniLutG31qMWYZ8PSI7WmN4E3Qnw
wJd2I5uRyFjhAGTRATpSZe1Cs2/MyDUlB0duJ8qXV7L9qsDT/L+P7tfRWfdEselfmMSfTi//BmhG
pk2/K3LJCBtxOTic5FJxgFSUnGdAndWKrvLPdD7NWmJ5CzseFMfrReDNDHLOzl3IsE6ZlWAKNi0S
kXb7P7UkGRthYPyATxuv4gzb5/1adl6QaJv2lVNSv9guzE+d97yaLCeBojI77YLAFioUKsZicLyl
huje4+/gGY79iCyWzZwRVSC4sFLfYuGWd2jraZfFQPBoqYKRdMZbHM5UnoQfGgYSIUdwoK/wD5rY
l/siPtP4gfTGt3eP6Rmu7LGx0i3BxSb24LqdF7k0M1bRmkTvjBrIoA7Ku+SCQoyPvPIAeawdmjwO
2daNGE7dE0NAxtvftpu5BUxYQxMOPZu0ag7dD7lMazlzklgbeamRlROP/S9XUh9mvN1Xi00CZtnx
TdryEmJ5qIOQrtVM6Ts75QVfSBnUqDbWa1kQnYPJox/LXZ/ngRhT+hJ++SWJ8ynKXCYQdPS4bf3w
PLC6UFF46If8lqhyZwFQWum/kLS+/F0CiUqwIMU1LtWHVfbsWqJnyu8zQFCn2icahLF96i5azYYo
mo7EI66I0kXVbAIOPcvdM56VuI+X9VbWKfTEwObm5fr7c2DK91yPNV3md+Kasnwj2GqMYoE1TbMN
X5GUd7EzuAJtJMlvkRHMrIa/liebbtdArezUMor8MfIK+yNoNyc3zXeZq0viy/wpU9HNHu8aQqDC
7gvoOoHkc/hmEAkrw827V68jYDVlw+Eb9pPPemt1/94jM1NQ4DxMr7IrLjYw1pQwrHSeJh4OBKXl
GdxpxYMMi8gPkBJyYyy7noloeNVMTE1NnWcNxVMhdUU1OCI6v81K8FM5edY5sWfER6HwcVHduy5R
LZ1dFRd0Yl/ya6So7xAqMUu+t/VpFVaLcjXQ83etsG0OaRM5f88EthmEnMfwPOQleoMMsQiw0fEa
CTOV0lDn2YP5+v4EFMmPrGtySiPnsSFLMaYxa8qeY3Keo57Z1zP84/GaFOx4kLtzikgYUlfCA+Iv
1R5C+/QbrD1GpSUIrmSDttZIiG10F0IpXtzK7ZAEpk2AiKncXIvSmkwtX1qa9AXCWEcc+B1gX3xY
YJt4Gx4XTUIGRJ3AbOZnjBtdIoMDaN6XF9M2SC9U0lR9nREueR4N/nPFIxBVgtXlVHpZ7BzbQrw+
Vee4CgJoM7rrLHwJT1c+wdVP8c/1d3HsIFk0YC55Cvudfn62+/BkBtjXKJgxqRQ4a222MKB98Maw
0TcGonvHrMhDfa0PHggIxMIQm2v+/4E3pdpQ7pxHbrUpSkzu2Eqiz7ONgI7UO/NK8vJQePC0oK0/
566K0285J9JLpHf2VjFdsmhtzQ7I2+LJT5VQIRJ6c4NfQ3+rr+mrqAikDtKOdpUH6rYgKfFCLdXK
eFqn96ez2g929awBOGanf78QA6qoiQUsYhh144qxY96d2ZYpY81788uBwHBWsU1flTtAKT4t6moT
bX3YHU7TONoaPgxDZDz7TfSdSgkHlq+nV+SeIlN4N2HJoxdPNMR6yT4pVVtGaEflwKzZiU4GzdQk
JUBZKwPtu785Q8tMM/5QZr572tRXDxxOQwolz763ckhLFJZOinFTm44nacbK2mkBNKOUORYDrJ/F
5Cz2SAeISxgkM2xpqpVD5kyxfUO8poe0RZDWQ4YDjy8/jrXyxbxclc4abNcA29vKSvg/7e6RQqy2
GOec7GJISkXprntHaYKLIg+2aypG5eWDooj0e4b/QUXrHqJG86h302MCkNUJRzzy9rJD8K/no7lx
+fqKeUgzU9bnrJrFGf++hT19rjYQdzN/nQJimrsOqeJQze+dAAud4GUMv7gQ61nsojFqOVEtriPg
ZAaeC+O81kBpATfrYhTDnB9GMegopvfGGb4ZLiq/yxVeN0ZCoKZHUrmiOp6QCfaroEdV5QUpdxcb
40lQOoyEH5ELjNOaH+Q5rFSe0kWzWNlMv3GhzZGBXu8/pwn8h9bYKmor8oQoQf69ixdZNJKhrWIh
Q/dRBTXiaFStFpHMw6mnmQrRaXyagEVXd+iXL8Hq2BjUPAUNpaVovmTIf8lg/hePFH3s8D8XRaG9
9EbXqDdc61rqXvE6e+9kgSdIt7nmhlz72GmvfAk4cgEIc5/YXhU5rp4La2/woHhUc/uzakflStxn
EL+b0orMzenXkKMb5O23dqAWC0GchY/wNADztY6x42WlZPoSDo3PYBUQhr6NAoNnCxIUECKddlqt
YqD5Mq8bylSKgiJusnuZxNxlJHV10iftZat3qHMKh5K46rhsQaPwqZd7SFp3mzko3ijLd0k/bey9
p5UWB92CDfBFRoL4i9v5kazPd3BMg7s0n7GsVfdFyqjvrPfY5Wnr2KfsHBdtfHd4W1rq/WdmhxZV
dxdC8LeP2xVKMdZAN+Pk/ygn5mkB0yAhyh/ZGvB5YsQPWyQhL6+2EWYt5Ne4aUqcEabQzX6Wh31L
lbFmS0H4ljsRq39Y0RLFQcci09uJZOpcjPX7n4KX/nM2TLYMIEnviu/BA92lAUXmCxrkZUh41fX5
v5awjaXVuelY7BG17H05UWyxnVfSuxO2EadLCEuWkU2xXkIsQPsaE8gAyD5qO9bLxXZ/fAeoeXTo
dXurJGIp+nUYZPXD2aL0Pm8tacOQS226LuY61d/hIZDKK6PMpKALeHFO/AvC2V+h4K40Ub55y/T+
ThlvwiwZhvloMuQY9FSzfmGZ7fDxUSbwI9TaaDp2lZ85MI56LmOfttYykyoYiVcUVKKeMHXHo8D1
XZstdO93of6f0tj6sv/qF/ws7xlGs1fpz1vlaxpfQwZW/jwMcK2p+WIXikiGnvfZnrV6Q4lRxcES
ArAEvMRRSJlhT9wrFX8m+2RV2nk45BlRVe/UTU29dqYHgRGhT61etdT7p2sbSrHcMEtga76FackO
/oEA6X12YZj1L7Q1yyJiSzMCfLj3Wtw09dsVJIZWSewbC+c9uRdC2L6BFGEF/VjyjdLh3pKI8krE
ufPgVdIotLc6fM6MjHuFB2k+HAwf0sIsYHn7udSOfSTVryfduE7olcwh6hubE/iSXBkClCTYTlJ9
12Nev1PgM1fRJigH3xyoa5ybN1H9ypCWStyhGJLbAmQIfWwjT43d651pc5blt3EP/wDk52nH2shY
eCpLkPanYTamzzG6g+uNAa2gr38BEHXKLk6BohamWgLCYBa1DOu2ouAXzDLykuBfU/c13oUCEzeO
43OxlN3BuokN53JPHxaNpv4F5SFlQgrPSo2/GE1wQvSk64wdyVkYbIs6cAC2NNt3ZXb9KSU232vj
Gb8TEZLnrPCRGaMPGN4SRog2gABc/C7PPzUIoIZJiZzYA0FnwsuXUQN7HWe5uDXADX60L4RTn+75
c5JEG2T5Az37V2q3XV9L62/KLBlyKvY6CDvaUI5xHSSqPSK1KnhYfp6x4ooV3wooltnGSTa8EteE
g9Mn77CvbOAbt55aroVRv3k8wdg4oqil8e/+KxMehACbxlWp0a1CtjbpLSJDcritkAOv7lSSKvKA
puMeOJyRfAgXwj7duvjrGpRJmikcN0osw2QW+gvIyZmFZwDh60b/9+5kIVlINjzyvrmnNVKFLRrJ
/+sLajnBcQ9pB8OXSHMXsTMQNdUMPUDsjmEWV7Y1zmI7HUOvv8NN2phxdvGzgWsbsICRqCXtfRML
FiJwh8BQdZE1opAdxE/i/FPZA032XNhnVaviSAeLv8BfZIm8gUE3MPCuMx6YsTVj5G4Irzvo11is
gLrAb9TVKjs9iaYy6tOl0xpNu0F3cOvCqr/j1uxn/MzhjtOI0rB8/1Ir2V5KRcN7m1iYhIgWJrCz
NE1JqzNB5ytu3PYBMcPavwen9NOBmdl9JSPzM28DuJJ//3vXNp2xEzi/+HkM3/f9mmOvOyd81aGD
MtiYhq0zlNfADe1jO+h5O8UjK8CBKllXCsfx3U+4KcQGmpmyObDT+YM0NXgrJ7Y/H8l5blWJfLrK
dqCBLKN896f0oOltI6irOGdsVbkcTQCwyH+3URRZtb45+WO5b/wSV4Zm0PKpq2Try5BvY596cbLh
gDkfY62TJyfDk4WDaU5vmWFuTcFr9HEB3MJQAcDnlp9QAwOlwjxz/hH//r8XBtAhoprMpxiarEQt
/0GpN9T4cIVH6zz9R6bucred5wHXUI1Lj6CjpMT5Xao8yK0l9UQA4IhHwPAOurEJx9qJxuYm8Zdq
zwRWnN3jVqTPb6ZUg+2MXBpOsN6Cx4hKjCXB7MzUN2RWJB47HhXJq6rOnDDsett09sm7djP7UnVq
wPHeLzwghZiB5k9RSJy4vFwfpK9c28kUqSHrpfUYYcZDpoInVHndN1ULvM8fMmoR1v8soGmDHBDr
OdZ7yYZ4ednaT3Vr785SJrwKmCwJBar5QCTLRyLJ3ZHTCvUrEz1tA4vRb2aYa8parnyZb22oxnDm
ZsscmbAo7OeXhLZ/D/7mIpOfiBdgvbQg4kvhLMRMqJBe+0FAmmJAn2bkWAxz11PhZtSlYze/qo42
vsa3NJDIXN3TbuKA1kflvKv3Vp2h4c7rgqVemu/QSKhfueiYPm+tHmH54jhYCOmghOr2APwW9wBS
cRZzqwn0o2fWtEgNo2gemt6R6rBQvpXlaJPvqEJhrtyL24V/KBAdCJ0fyEccaos+IJ9JK3REL0OZ
LCjAnzhIIa9k0t7QNiFJs1KsqpMM7s1pteAYAC+rpKACxZ8AQSBUQ0y/C4hrIj9JDL2ZxGriBVHC
nYQHv5tLsQM/qYbctsEI5j3AcCMS3bZ0jD53PO5EgoaKQJ5BkxP5FKcjVRdStof92wkKq5v0SrDP
HKr8epgvEzgnG3EgjGCmdTnEQZESio0VA7zijIqLJZbfAu7XP7co22F53WdUloSUcpY0NChoMRhl
JPFDIxXOtC2ltYu6QEZ6DtSvMKjk3D/gJkVpiJiBRGUlbmdzxDinmtz298G7BP/YApmdmUCA8jdN
tpmFAlOCTVlfVNqEX3ADanfl4vEPQ357vcakGUX1Bh1W+eHFiDRZmGMdbUIJr8QZuoNqkVPFIonx
lB3ngf6ovMKKhKLoAbcsF/mGfW5Ha8vj5yaaFRa1O5batNxCuvPX31U8iWO5n+oChwFQbQD9wDI7
qHGgwiMAEP6miLCI/Rw8YTFEWQaqaH1KY1uOwpHXk8j28iMRVn5PaVikHeG7ajUJY1LnQgBWq79w
BP0k6cMWr/UIMLUjDPXYnpxEmQdRYLUmLDljARZcGkf5Qr7G04klH8sifIF/wH6sVlBaTOSWHWLX
EFG4NfuIgC8jsTwFnEoxxbiwwQ82MH2wEeYuxxcG6i8/KGlLvjTQA4uqU98XYXr+S4TqhcZWCixi
Psnl8iEW4et2+A8DsQvRqxUkzhP0DDS9RSXH1xefvu4BrnJbBBaLwulNA5OnLn6LBAnNXGSx4MyS
69XSc/WTs7Z8EVuxTMqMi8Huf7wf5PTT1vvL5Q7legC8j/ExQpmrthOBivnq7sX36CoRWx1QuRTB
xBZztNaVfHHz7oR5vChIybiJ+LjGXuOw89qK+Gz6xir2mK32LKsPCbTvt81q4TKV6qNIy5/ME+Ad
jU/gzIXGd4yoTXLKviWICWhDiZi8tUlo9mzeU9HLb77ue0xmfhLTae8+l7EdmTFopnTL9Wl5uUQh
YRQsYB0ygV1zpPrZZEsjJ7TdZKDCvVZ4F698mkvTnEF6bawqbdyQm+7EZnCH1njU03+/IEYQHP0L
MjZgXhFM+3dtifHpl3Bj1KdpI+O7AAlFp+gq1DUmsD9E3aAKgOOoJvpjYcJ9f6tCFL1c0+ke66fD
snZfSAr5lOjQA1hbcI/tAzMMTpqglQWjs1XyKhQKvhzDZZ93kB7wwP9K0XG7K+5T92Dn+57TiHgS
1InNepJkHjhk6D71k+xHZoioXSh9adQGuFfrt5TF6NBAXZmerM5UEtU5UiY/TMyxZ/E5LgKZA1Dl
xm1xrBxRbpaIYo1LAPKsR2PG2+pGzEdoDmqtNQkN7sTDUKU+GFDvOs7ix4hmQXxRcugCUOO0R4Ig
H6N7dqcBsb8iu2oc/c9yu4mF1VneS+6VkVJt+q5Ak+fv4Z1LAApgv1J+eN3PZMeIc3X0ICp+OGw+
S3HF4gjAmmaQV3UrbZipUIFmcP01U9tiVpa6Pru2udyC6LnZ6Nz06PM0wAgNCdDcWsOaFOnLsNwk
ECst+T1VOFMNGpxzpFAc4q11ECir+bB0LYGT64vkwdGf7jLpB+vhSGKcYA/E5HI064Bw7sOM4/MY
Nu88t1Rk/Lz+tSpP7uoK2aRz4XAXdVh968RFfh5JwDie9cFXElS58oRoth4ULKWEyxvyIGkXfoXw
dfpqlTJWNx7LnxCVT5ulfOd0g6xkeU15vUdDdH3b3FkRJQFhqgMXMFBVnF2moNHNxk+oTBbs2EtM
P6qD8mwgDv5qKBNCWn+BIHvPQrKT7yQCW6WNzxjH/JcbuBNXwWkMkUCuvXrFIZW2/sdeAvj174jx
S06mxYQ2Vu7+J1nPXJA11vBH3GUtLg0c1ddd/+ukmaFdao1v+w2c/bEmsoQSsv3THB2RFD18oFJS
O1XvuGIjc6g2PvjD9Ea/yTpR71lIAQxefAxHnpnckqFz95NsxDtp/HrzKZwHb9fCDQ3Od28lHcp8
LMLxDnEFwjveHVxZMx+sb2PnoMJYwodcKlWEcwfqDX8fKeAvKQ+fpQNsN7MZnCSbJInPXosw5y4w
IVQL/HIni2sqGWXqm8OohDUn35UUTL8sLqoDVJ/MstLFOpk8gNxxS+xS1GM5G0/+bpQzcTRppKZU
okb0BAdTu14JLeDppGd20y/7/lHRrM+L8IRGCZ+5UBysXi+xjT9V3Lk82G5CJlYbeB7Lsi+Tc+lQ
2JMycyTvPhSVAw2VyxM+BqmF5KaA8TEbxWKqZul2vcVoGRMnRi+6MDjtKNP2IUCY6Q0+CRBMOHTh
bmcjQ+IOoR+wULe1Z6iwjOHj6fUP44W18p2Cwi6OFRXeqc5fBxtBWt0YeRhfLP8Qs/sVCMYERQZe
RjijYH+iTHVTsrTnGo4kNq7pRbEr3fzd85RgtTX18jJRSWyuyyziazTOMK5EIiT7LRKsEp5NxSMJ
8O8clup/Zjqh2ThQoe4paB4HgoxDp1GKoNNC82Ys8Fbn9mr/R+3PEGyMsdGnIgL1d9R3zH93PNgr
EE2AkwhFbOE7VGPafIAlFHi7Z4pNeYvta0ycZHXhuWBLJsPkXnYFnmS+S4FPMw9YMoeT+ZCUPZJd
l/YSneDaw+xiQ2Bz32n4SB202x3iwx41PGGN/n/njA5wg1xhSzSWuI5+kt71lCfvKNFMJa4rm9BM
PxMMMy+tDBB3opaN5g3balb9M59n0lF1HdOnN+bUndacgbJap8pyekNKz4Iouyy1H3YOtzqLW0j5
ksaJS7XQaOsZklbVVBi2vjT3Qldu+TqjQz04mQ3E2uO9dFaYgqRfapOF0IxCkQGJrwmiVYW3pVfD
BkoE+LSxBZG/fYOipsPvrRlkvwt3CD7eD9ixl8VHkPxXYi+/sFOFIY5aW3g/9h+mt+rBX9BfQ0n7
Szf4vUXYZmynOk6Yxkkb29lZ1V3SoaujGhgBbsKJoItdpWMcWZdcSEj5TcdJ9sP7o5Mw2dysf8eU
vJzOEztB+RR+CKCv4jjN9jF3wQS5tsyskzkuh1f1n+xbSCCmByoArbMP8vh0e2GmwhMsjYj1tkNI
d6bk49E9PuRpJVfgPDvMNQ27AJWds6BO4yxzp9gqkBm+LnB4Q5YhKnQWPcseiqL3O8jf3BpIpFo3
2g4PZ/7BzECqyG+pb23PDlNRBIjkVsmQzPLTqfhxvv9P3RKufVnM+pU27YTKDpIrcptfP7z1+iq1
JbnS1Z0zp6t1VGJi0z6oJ0ZlY3m4BE14RxmnR7w/xjh2oxVvUoIyI1yl9CtXLwO3AHhCzQGLfivv
r5O0Q8ZC/3Z62aTN4/7JvwSqcDm3z7dc+MMe74N2pjjitMhPYQPjh8j7jH9tI7WqRC4NhBJsInah
AeZyadKmX/hjKW3o8kLrlbKOIj/cyrvRk+Ij3R56o2NXv4RAIizMmPVUSTsA2xfo9YBLYYcNs+6y
B7c4oYpM8vPcL2fOtPp6nrietzdITEPULxaGqVs0INNxuYJkg++ew7qWZE3dtgJqCmSXYc9LopzV
eOe6WFiNUuMTS7bhrKoASaSLXry+E778RtacMFUyRxepg/yrIIoDm0ZUIMYBFqtYs/8BWGM3tDDI
dqb3x5XruRdfVP724lo5fzg58WoNe6suBvIts7BmZNbAIDnohkMjwAYEXinVvTk55WTFH+EJQSgO
uRM9Mb5aY1jgzD4y+XtThovK9YFPiKh5zjdDKyGyRto0aUiTviTsvKDj+HdRjIhERKQREWgFSrGm
qZGlT6vdpzp4rgAzt4IOH4r60be5nQ/STDMdfCG6IQm22pn2YRahDFcrF/Sl4W7SdermwxIeazj7
hKaCT6rlsWrOgwdgj0Neml71SSyLpr3hlBRs0XGjPvnJPN5KeT6kTiJ4xC7tW2+iaVIXGXu00TYW
oErChM03m8Vrkyvcch5ZQNhHdSCzVLLrmF0HU1VEDg45V3iyxbth0PK2vChflCL/IV1/5UakodTu
lnI66kXZFQmhfZchBTCFLI1lNGTgdOlpTULIEZfbee3FKtqIFM6daox7ppJ4Q6vjIOq39QukIyGX
RuJDsi8leF5/YLS63uSAEYpmmhYyEoLJ1/Ngb901OkPgr9TPQ5q22JHC4iBJgFLqRvI23tp7o9ba
AjqGR1N8OGW8ksdApuAKQF/NDhuT98gVw/jSkW6YRZGTbgPygNPrAnabDdo/dxMN8So8kOQ9lXyY
ckXFrT6FD7N56GAU2z5g97JtTv/rR44l61n9KhQb6PORV7rpvj37sWmthZep98ZiQ5cpwFBYRVBa
/2MJklO/TKDoMkR0YKzgD8au+hvR7Ot7EXswS+Ay9THcmbsPs1tf37WcIvird3lQslhGptqgj7UZ
FkFfwsKlFuvZ6qC5Zqvd01rmH7cqMl/qUr9IxUYE0cVh0XE9R3MeYoQuxBLKjNOEDfr6z+lGtb0W
EcJFq4iln/lSWXcH4aS8V4ZQ/BCKdCNuZdNbF8VXeNhDIIWwoq6sKuZ8Glw/XXuGQ5yGGjDxWPQU
x/kUPyCDh8MCs8bceb6kn+eY0zDQOdAh9xuCmSYNJ3QVIT5t5rXbm+y6GKV1pDdipw6dYYsonl3Z
P95x1FvBTkTqVCUJqpKeRfe0ungV1V8PPV1w82dYJq5xp5h0jMgfcLLQuQKyhxlLB/HaKGlzC9VO
6jITpYB/BRuPmr+liZr9tR+QTQKPhkbNdcltZ+B/a0tiQTY+/ijIN2mUAgGyrYlguMcfomXPas+T
kSTQU+uCofKNvggWnWVXZ8/AR+61LCtfdVU1MctY16P2Ma7YMx+iPvfKXj1LZPw8qVnch+kENzWt
I3mByVyduub5hRFtYr2CcqkfMBY2WQkdR7cwBCav3lKR4bPk5oEEHqusOzvJrrDAwlO/Ev+cJU3H
8SUr5gRVNZSAUxXz1ec0pszMe3ci3mnqCLu8MHIu5QHYb4c2/1QH58r/EB+e8up1LZAowUhsazKo
t7i5tJRRVM580Sn/GkAZrD7bdh/dWN0nwQNwl4xL/Eg6RpBk8cteowhGAeYpnq3O76+jPmDOpb7q
UWiNVlO/tzMHK905AyxUHntVYJVC940K+wdpUB7IRKP2YVmil9W6gN7KwZULei5iRxke53zPdpve
LqV7yy4dg1nZyZlbfZ6efHy2BSzFccxPHKcQxQCDEOIfsdNPyt1WscJufelKT8wQYNXNKvcgpXul
ZC86sFKx8YKVQYaZieIUvIdT5/i7slEFynWfQWZaFblaCMu/VL+szSiD3FEWXcBnIkYGsoc3D14m
dNtf4aLRI1aLF7MJSjqbalS4IBp3NdI+JkTKTpHkZg7LU1Ka2qXfgww4ia0575+H+BQ4UnhnQki3
l4fb8RVxN7s0RTTq4HQv8lqg17ah2w925ys1dpiCUpGusA0YD9pLF9/eKL56sqSLWily4mRW25lY
3u/Awk9lMyv3XECZZsS9f9PLkndqZaa78QRYqFvfwkDz/IpOhUYTxsISHmKkmYW/EJP9n7CPawjH
VC3ldb9G/rFxLM3mDN9rs/xcrrLlcEMaBcWUSYdL76GtU93tr0S0HlVZXoChPQweNPOlFm0ZHl6j
RJMgWzGeh8dCbI00SfNUbdlwnK0P+Z5v6KEFCjBKZny/ng5mzJVS1yEuKhXEos7dEbtUOzOlQL0c
7uvpZEw62khZzSK6c7F8HAbCuUm2lXUGRKb1OuxvhJ7ZPosR2dOKOGphivOnKOmK6g4cZWYX6VnF
J8kzqT5UTcZ551I3jnWbgpQiCa1eHIV5ADqK6+zhS7/rXfY7tQhCqBWo8J+GBEQMhUMiPLv170xK
oj2mpqFkW4sgZ1/MMMHUAxtoy26FCgf88XSki1qwrw9Eyv5h4W8Q48mbuj24aIBfusrRKoH1b6AX
PRHlHjAkeRDKUSl4OkSwao37ct2hQ7L2sji2ahy5hbPFu4Kw2P/lbSp8L+KoxWszHzueSz1D4Uam
tWPFNPz693Ql3KMdQrPjOrz6DnleNM0N9hy8CAdi+T/jtXQOu7xg8b2S4dMY8hMB9Yb8aeoYbrnZ
ZviGaUnLDX0wVjMd5R8IXqtis2m2gQCDhGW6RjA0AG9ldhhHZcgrAMaFwGFP/agiHzWkeWDPb45d
dx7o/AoxOE8suAlgTMnSoB6Hw6kuCKLb/rjyemYMFyy14QTv5Cy3nFtE2bExjr7CLXOaDS1dKSMf
dGhHBmswQtE8VW9nR8v43Tp6m5vocUa2d9uZ1IYvjp1Cz2RwsV/h1aunuDtAZZi0sWPQ0r+zhmGb
2LhNWId3g+jIW1fbThYRQwLQMh3E5O4QjY8D2W5FJ8cmEYqnc8vu4Fz/xQ9vbELlK4NYdQU9CBnh
8gqM/o6DP2HG//GfjTdHQfJ87bemwoamgbVcEQdvsHVoEgO2NfGHpsc/2g0AUwfgVDVWMtLRMLVX
THY8ZPOHomEoBG7a7Q+JGEhvmgDUz+zsshek49LVuFnu7rfcJAB18YTxqFU5PD7B+b+NBqGaBRBk
XVnhU9pWcMLWfImMYGA8l2xgSL9hWDAO9ZA2zCPFXFika0OFUFbMjIlwIjce426qUV3CgUvDCKCN
O7doWUAyrMBP29Cy6Uw1gFYi5VfiD5FxdU42xRx0MuDm/Orf3LmCapLVSMWwDLuIcM95gfTd/pv/
NniQAfScjEhAbbWZ+3eHA+j1/3qnn5fD5sQyVF9zVc1Cb69fA4p72Q+s8xm8QJWD9rmUAip0UJ/A
Gs78SiIXNdiIUjsLrza1Ejp4AXfwbiraqzZ5lyvOJiToNvafMsne9zQu5Pny2xPC0Hgu35nIHiAd
waLJeYdZ/PKwUpmVlh2TSCzDGehkUI1xS1Q8rWm08SbKM5b5G/Ea9Om96M0qfNSYciLgnxFzT82t
zyuV8C/2Tbg+DTwXaeIEWc3rvSNo6ZqA7C/2zHwyMq/OKwrLLExSqiJ6nwi0CkX9kTBvtAm/AOVc
QJ3fKAPy4S0IAvSH/2ozvble300FIXc3OecvywUbNqLSgswIsSyD4BSM7Pv0ekWZWR8O3MfoIuKe
U8yUcTIttn+2ovCMsxf9nAldEFc/md9QgFcTPXKufnJPrBpbZMzgLdfoXDS7bOnZHgClSZLxGBrC
jFXBmX0/gKds1qdJT7UOVFEWW7ySpA6CoR/lS24zY/W9a5y+8H8YYNpBun7OeOgChtYn/XZOXOZM
+uws0uWTaLurshIIUYFm3S63sa05aWbJv8dVgCwD02L4+cA7E2sd/roOxSQ7vVkCgx8fi9+SCE/3
Ew+lKwEi93No/TQJ+XJcjymXsQ/T43bK4uGuMji0NtGnw2alrgJU/h6CCDn4j3Oq83dmpGuOi54T
/BxwD1TpfAqiAiwaMLJmGNh9NPrqQCUJo9NWub5VUzIspLZUPf6MaxZjaa6wUdN3XmIYfMVXy/lc
G+NKiYVMwhB6VSb60Kt/wvibVE098LhQRzqjh7fnNjrAE0BE4z00/3l2dhrltnwqD5KDuyDClxqN
KZMiNiu5XKq/SlHcl+xv1B9sbFoh7aCSxDw8CoVxUNFpP8La91L6uohgGrcNQvuNpd8OftaX/ym9
08Y6RR9xGs5j/yJ7mKVB/yJXGYNuQ7d1n4H6R3DIM+07wk0Uh29BqH5IX1vfIFPRy+cgVjm0XBmf
yjuVy0NGi5QsaF1LAsBDbAKfaF6QFFCZYVcN+lDtNCHCsRvFAWPH5d4/63GSw+P5tXH7Goyi4PYn
710gdeClmnedFcts4hpOg1CW/gWt9Yj/Zwg1kE6O8LoNjifurjQ/Gz7Uwp47OGXteyK++2IyrWjx
aLX7JfgebhSbSXHPH8bbxu2MLKcNvlL2+GYa+nqZphTr65GI3HSgujJ+S6/G1UpVlBkJLsAdaPVo
ozWdv721+4sDmqGduOA9s/d4wwUI/RaJUZZ2HQ2XH265uVNcSBpRYw+KbPhfPp9LYJKcQiVd99KZ
ufvxMU9acCaSDnwgVJlVhoh+11hrXMJrVLn63k0ddW2e9Z2TD118SQEguW7bQpGrN3Rtzo9HSubz
9BMos/ZbBpBI0h5qaTMeKGiqgRLWOeK4332UVb76OxneRqiFOXlwUy53QGfNU6RsqjqFKt+Qu1tY
X/LjGhXsGL7YQ7rS+qjc9Q6oaXTnJoV8O0S7N01YiMWwJ2phbXqCJd56Pnx3j1mgRkV3Q6NcmHgB
gUqfGHqWpKz6E29Eg2m0TrhAW7TX+jTzpbECQMcmRKunSbUHTc9v1zDxL7FLsCNpKoK5HEveW/c7
y7G9tjBXIA9oVv6/LINxUMEuaLicwgGzSCmjNyev2jUuZvDsH5Rr3U2OjFBcjbtzO8dGw37kKIv0
oe9JHK2iTu6j9vo4tGqGYc9rw4wDss11n7Pr2NFNTxlXfI7OQT4ajAiJCAT9KGBuXahg9xsNR/wt
+D600buiGc+JsSCZJmuu6Jk7CdgPKXrooIIc/dU8RIWMRxPJQu7L9ZgXkscLgEF93eWxarn40Tfp
WWV4+9ULbARI5Sjwe9rAeOfqqZ/A9i9vsjkwUFf9LAjSu5ElteUy5+ISV9GaWDmTDYMbNxYrI9Ix
YiQZiPXeIHPo/1z0wp/yFMPHlsLs7pBTBzKEvxthoAP6SZUto0ydin+2DzRjJO4WQT/1WXTjmWnV
P8MvVRLgcUxLcCd6I8BkXYQgqBfC/b261o74XjUUjs2xHiWKe3XOQGa9Dhiivzm34gGHzYGfO8zB
CRDTEFOogmqiDrHPBw2ggNyufFNqN0Gz90y5LC7GIhediox2geQ3pwzGKXZGfO16Q7R/EXkh8A4x
ffkDMPPK2PU2sT62Oni5y74yq+Z62ggbL3GkT4L3kpNjDmq4QHpXnB49CdKrpJby1idCFoMJa5JY
K9vUK8NibD+QYU8N7HzRRC/zbZ5zDOOZfA5OmDbyH4txK6qTxC2cu6ojom+qGl0PQNohniZmNYOg
locAnk46HgNyokvV1FuYtFH3x5vR5QXnB162RAjz66rqZiUjocOlb4dW3yLCvMG4OtG7Z15zETaX
aJPFCtqrfaq9rhePtfkNpALZ9f7fz+1aYyuVgqZo8kk9vU2znLYW2gpCvcCGta4wZlHrJWOmXH3o
0CkgYjlWQe8D2p/4vtBvCW1+PdNPM/mK267VsNXKhoMqRzK8faozP3HBQoVGBpdtIkO6CUu4QNBo
h3NoBLvNiVvrep4naJ46JmUvqzTmoh6+PXNA5jbmdJuf0vZt9k09YYghpvqHZu3RSkca2kz8mZHq
GncUQAcwuXnCnNgwaNR9s2tYdAMTURZmLqtfb657+7TSBwzQHbT0WzoJGiB3pJoPCl6wtKz4y3RO
ZwRY4JeGsCOcXq4qYlSdpgDmnAsg5tP76ci8K3VJaP2X81Z2ZuqEIbEeLNfzrXcq/X7hLq/FN6ka
HOWsYI3bIH/80DKT2jtPHWBQuZfgiOLKBNW52TNrCDwj5QYSdivq8rXa14A/Em/jtp11BRZS5zBf
mBKcj8tqc8k5ukKUzg9YTTBtVsVN5lEom2B28kAe3s1bQMILCt1bNwY9yDWtWCvNwGMrBv/XrEXE
wfxvSHksUxqPaA/70nLOhh3Sv96OaqjEp/CHxYJk2/er39IRBtUpO7zJjrVj2YogVzCRAhLIXmcE
pdZVxXzOl4NSuh2W3UEJgjYirq3FDiyGsbKCIT/Q3Z9Y4kzDj35Ln/mIj1c2RsBhQDohBBELeSwM
PYzRkTfGJXnXiBsvpgoGND+310Fii0LK+v2uJjMkX1kSNKo8y7/uE3LCgsY2B2i5xKUflwkvK24w
2SevPGPEJVr06Os9Yxfp3nVinXHwmoDLQ+h3zS+Uuy/JXqPah9YKCS+AphU/2GNWJTgIZXMru2Wf
wGiEhBwQeOtBdORFLnwaE+loC0LmAjFyvaUDYbCkgy45wzdaup+y1qj+sMNbe7SUXuGOQWGKoJHJ
bj/LSZYBu2fbnxyxU0Okfb+mFeytQ7DhYFC9ASMWFJXTxJkA4GYHod0vnZjzV+IOxyRJs9tasfbS
etGw9Xs76fjmIPr4oP2MxmtCZM0/Rq7xiJM7ZN9l9Mdbm6z0YMX8s38EZeQPq8c69UjJwDuYsi7y
4n4ZUxkgp1IlHw1ZHz/sJOD+l2nFHsOZlQZ0XKcQhcR/UPjE2XwKnNSJHdpyr1qTD9elPVq34/2l
Gh4kfir5i59vvZwB2vtt2i0wYkaUB/jWVSFjbmNteon9x4fWLFrZH8db5930ZCsyJibSmaCfi9h7
w7ciEVQgDYhw1vACINRZ/MP5wZVb7yc4dZPx6st9ce9QZsgH/8Vp2UUDvPuomvRjDxtPeoqw+HBW
ThbHEv6zsrXpOJCj8hYCChjwPf+WCoW6HbxD/+jKSD9OxUbmWmXg1E6UyT1glzShCIFGJt5EmxPk
ykBwZRTW4rJ06aicXRFb6dfvCknmxvn1FrDQb4ih7XYKqCEqYs79h0l6q44e3w2CeSEB47/ZvKUc
PcJ3uAWiBhgJvpaGJ2M6eGIfnJS6bfzI2OCGP7kbASh4Y66JOCRGiKC1OOben1zbxxneh9Zijncx
mK6/5vyVXK3xQysPIS8H3SsPxI7QZxvBAzPgliAWjwm2icST4E6qdfNWXAxwOcpElLkuVQ1fmO3O
0glob8yzGkYpkNg8rFx08aYbu57re8hX0TqYh0h11aSdPo9GPN+v4PmxSxIb3AcY0lEXwjX8SCmC
GYxSrToPDXzxgo5S58ejD+Wf8gZspx6wd18ElEOApTcqMYN54EyXZOE2BSKqsE4C6Ff1I6gumECB
o9aihkMjlsqI/Skg/uu6uaW4/Nhq8p6fna0pAAiLddCgzAmZ8Q9modG4StNyWDjh0lxBEZPZQphJ
Jx/+yg96jFOppZ4yPg5cfTuBrXVwBDbmUOGwGBv+upUcrG7nuOVX0hGjHhG1SwUdNDn+G73XNiyC
+oyIsi8ff0zo4nYP1pDqeqh+QKslF7lsbCEDz7RS5JcCZEhhRiGOuM6nboXvhNIT6K7mfsJQemmX
MvZkO8OSUkx6+4WuIfQOE2r5sBCxTv50v1Ke5wFgvwPlcYVTPNpENr5xxy3CNM4eBhNrhqbT2DpI
g3kBvUleuKbHzU6hJ50o3zrFFowd6FPKXCLSILT22bUPgSGSDinBFokeuhMXrf0pjRWe+gEpWsaV
9TNrGY6avtoiuKFnrEy0gdkW/r9s4wZU9wuPpbG2mNeMAVNpGN4CXoldl3uSwLwQnLPTp7eIRczm
VEjffW1m3sT6SOmrpG/iBATeAt7pnBKGKHiFTFkW6GSFSyQjP7juDX5snEP0JUzpZ81nsh7Exubr
kWk83D/MZLKpyzxd2RZ5YzSDjSL84t0aSofpOsoDm8wZZc8e9eZIgL0TtBTMnQ+gUDBSmBzGPGjS
BwDMJgpADhRxsStPEErxy70lPjwi2bCC2N5WmY6+0PqXivxkubDrqxDnko9tlwaF+nPNp+4zjrRj
qTUogoUVUnlsPfRlSqpZ2AzxLDbz2mwdeaQ0rhg9HBjZesm1v4PFpEAAll/wlhQYfOM3f90dFo6L
6/CWNgsTeO6Ce1+JBk3zkcVgUVUlnTRpRkRPw9LvdNcHNqouyoX7DxMaz5km6wcPV/ft/QBviD2g
P8XWkSrCOhT/obpX919UXx1eR+iGLQBxDOINwVeejVvBj2YX8jNMj5HrwmoKPH0ZmQ6H1qC9aTJX
OLI2KfAhXSoISoIEmWxQMhrrbaNSP25n1Sn0S8VKUEeGTiBO8P1BF0sbtOxf2Tgz9x4ZbTGHm0YK
Kw0xjQINssJDxu/QeEbxW6W0nPMLKiH/QTd18CRSsRE/Jj96WOGBI3ScthBFzsVL8tzc6zfZv6z0
hHDjrcycnVayk428xgI4FdTqeur4uKAipfP5kpHExi1L0oxWHYaTLPxiDRcwq8ztsyy+YkNtdIsg
UjH36jl5+sIU5aIlcYjBAPDpVDIx3/LdRLuqmoKNGr6JtuaCIhdJ+/qyPLXFI54Fex4WTDNL3D40
ipbg7Wx5KhvLiJn9MXiQ1s0tZD7i2iJ6/qTzZmXftrm1PtNTGjZ7IHPKRIlFhgh1ENv2xc7UaDYG
6zev0Nf/WbfYxs8tTV3tKi3VVC1pri6Qt5Vl0ox4+OVh12WpBn54TlbJQtS7BK7X6q7zLHa/pk+A
R1OVEyJQ/2Vyx3O2+OxFSWJa36jVLbZensFnC5HXa8nfxnJrxdVnQCbvw4dLMAIl/zvQN/K5hHBP
akn81XkYx0d2XWdkBQeB1BjYE3fSy+j6Qv12oyFshwFDjrt9O+j7XG+wowBwCEzbdeZXPz/CtnMS
DbmXyJHI4Bc+fDFx81wnFfjooOjlqNuj7IN8Y6dUW8p6VlN7rftkCAg5eA7NezoQFVABHCEqckKE
8uPoxCS0VqdbDMuDMoh0L+FWZhMVjgspnTY0dgF8zrilw4+PKq3k5+3Qzm10xqT+O6L0izGGTbC9
bcEuwQhQvI5yMc/8k11PcJMjWjdgfI6gO9VLO4f4SOVTECV+BZOM8DE3D26FQqnCisNOlsToAL7g
jwZPBgIRZC5eOB1fP7I7Kr59J5z9p3K7aRw+NsrlPcu1IgJHm5zfx883vbDm36qdWdmiGq6ywdkl
w2mcBEbb99iWBE8PPTSKF6oXsVzyHwnApYcaod94MMaNHxzWa1mLQ/yrvP+23WCEWdCyeC5Xlyri
43t1SSRMgj+YWHqP2MShlK6cHVhXeuWAbfbaml3uaETMgRcKewR3XNmCU6ICE/kKZMSRsllRdd+M
OEiS8irSOGCl9Gc21EzBQkc9WX32W9phd3uReWGsG+ZdVs7di20WySm6yLP/tBn/YP6nDOur+UIX
+6Qaw81+/9gFvfEiTsBdXslDGQC9nnNUbFwNy32UwhMZbdx+OeKLA0szsC0qoXKcyMwlCRncmVS2
04djd3OcP+nHwKA/FfaXVozFTI6IX9fUXDHkkziO9h3pQ3pXS64ENeCEO4PfCyBT+3hzllUTiFJC
/Om2yDTth3KBeR+sDUaGdu119SfJ5pxgI7DzL/lIn66fetgQ75chEloaESoSFL5tiokcQQrLP2Dx
qiWWxmZFAFrH1raZcKcbSl36cBBtumPK/O58neHlpHX5Ot5ILv+Tx9pZJhjSpBdeQNbXsbClxpsI
tuuXwRkMYHrKW2pGNwicrkrXCgjIfa+fYtR5YoR4YWLy2hYjuLx68wor2UNvDSEU3oxHcxHDsvl4
9iL2VUz2c+Psxg6UWeHwrll7ulLouwBGBseqy1irHaqu7atKFz8GOblfTkdxgbOdXDuAc+PzftEE
Ny091grtwO0Exd2CSR+kyWwTdJQ06N9I9GBsIcGLk97adDYDOGSKcRukyA9L0I3UxT9Z1tRSFNr3
r96GkHI66LeWTKnzy9m9xRNSZPYklvcr27infCVoXWRTnLSfSHzPqHGqF64mdV5avoPtrgrDQ3fT
4bfz7AJxpQLxmxBBoZe46UVW3Vq9gvoIUwktQzt+aNf5lrR8/zK44bDRfh9JVLJh2L7N1EYAxQWN
AlF+JAcnHsPPBpU+ck5LqZwiXQsQ1uf4M76/y/kYKtNTZcFRrYCs7Eqdmu0J/Vey6QoiJWuozliw
0QEqwrFOUFaV6Eto9/3AKY5kh+rSoaH+pLB7c8IGO8jLexaqa5w2Ht0T8xEs//TcnnMT7aFQkxs+
TUcC1PNx+beYiDYb1x6qurCJdzGASX8m7580Km8+JuKsXLCQkuaAXEpHLw7vSx/U9i5XrRQtUE5r
Q1diODRFBN8eGud01NuhjvUtqHG9KsDiYsGybQm5wks1Si8LecOtdDDWWbx9TbL+cBjfYukSxnRG
zsV65RxGcr4jbZ3xG8l+KsGQKXGh0ldVvFOmZTa/WulADuSoEe8lOQZDGuLAlrhXHCmSKaKDcpnI
dsGgZbhOGLzmLjIvxPDlKLqGUGLpvGoNDY3k5+vN2e+Yhpc2YxuyEyIyne97rjCooFDoXN0QS2Gk
T9AA3v1XQphzCn88L99UeCNDl8jxl0+YPqc/Qa8OUZHWQw+tnMtSy5w5USszlu6V52mmvVJ/xFre
iMraZQNGmeVR+CmlnY4Kvh+eKoR8x7NepWeVaTMUjIku6cGBlvmLFbVNTZlQeiJ5hvROjTfqbBY4
F6JKOUEBqxknIGUCvyPTDzkySld6x5l2uf5BBNWzAqL8gqTL2wPRKZ3m4R0/ZtMPHO7LNI+2h8io
LTjpFng2dkLFxa1+iF1FhMZBr+KBFa1ld+rDloXyNVJATi4Va5oLhHjO03yy72sW4WNNZ5Jjq6Uq
e6FTZmI4vm7xasD94upBbhzpWwFrpoovuSofz1eMv9xw2enS1cD3eGsCMKyVYf7UZAitukscwKYl
bLa55Z+gNTmsp33WK7qfp1+oKGqo9rsP4S/+rEMHgFHheXW0hXzirCmlepnYrhhr4DFPJi+AUAhh
/rzzZVTbBO+07kpw5Hq15MgSa+m2b8OKW0ESdg3Wb/iPrWmeyhUfOQL8lP+gSkJjXV/H15yCym6Z
uBQBQiFT/2xj+2VYy0Nlk6jNOgZbpZ5MkEtrqeBvvHV7y+TuzNVlWgVWezT9lCKW2aOBXO4EXWWx
WGM6i7Fp8+6fWIJaTnKblnLCFFtGONjdMk5jq8h1vgODsPmOt0VOSZMAvAej4YvYVERQYiQ2Zqgz
6NWQd7c8xj9Z7QOLJBv8X+O5rx9X8SNyWtIAFTC1upcwYrjKAobs+mh9CwiJMkKXCfLcnuDN9FLt
Q4ugq82Jo+ezhs2yaF5lORZntWLgSLdqRUUNF8Jvo+0pM31PSFoLKUJreqsj41hjrWJDr/TZa6rQ
mUWJxmH7AmuMwkcuyVVQE8IHv/Oe1ay7N7nXOdgpXYrmPjtwtuGtiK9osRnMmC0GmRpGq0RsTQxA
QtELDTt4MXKLV42EXqv/S3JCK8CVTqG3MYqiIXz/XlXwpQSvwIGd39slXVHtvtpPJYGxUXkDUFLA
LLazPUhjm1XaxuYkMRDjxnt5AJy1Lw7SvJHR7ykdFhn/opmDUHEFiQVJlkA4HIZlfXgG27ZdFVo3
ZXmKcoshISqpPCFMDQMXOdLsYrLjd5qrb+5ZsIFEb/ES1PNmD6LkXFs+r9yIALCZ90Zq8cB3XPMB
KnoPR/RinEz/ws6DW4PNmifREvqVQTMd/Sai6rCchrONER/511tfxC6htCTiKCzfNmBgAi9iP7Y/
sJ7d7GN7afMzcjyGVxiJ6IPXfbGmtJuJw4KX9bzAGKunM3un8cFpr7poOi4wWB6hgAiu+jH4ftMr
ZAgxz9UQFReE2fvIibjqcK2wB2Qz5PA4LOB9G+kQqGdk992ycfuZAvnpxQf4qtxws/aqf1k10+8B
uadaH8MW6v8o5fDWEP1PNvdkhyj6VqVatZY4JVdHSPJitW221hq+uAfn8IXR7AZEmcvS5D1S2IdV
8zyDTejwnRF/oLc387aD55ehiAU6Bix/5QIitOqzHzx89Rr0JePkvS5qwodpv3ZvUY5MqnYU8OjN
2p1m7YXUAKdWmWZtD79RdZZrskpE+XmV0SgYIFUR2rBw2Mro2xzn+BToe1hgVzelXaeT5PLJV3VB
1h5Q1CSDBCO4r/3bsa/JEOWXwBFOhe8d5CHYW0eqNHZTP6ohyXrU33XsLMbtAbtMdvyYQHswFrF5
HrD6CUR1Z2k/n4W6yJdYWPPCF4nTm2qC6J/N+/HvoBU6UqcEtcESTxQgpz/DdLvqbjE9HvFTzDR9
4cJQ1QMWV4kX8BLalk/BzzSdFQ9WqP/ESpaxEGgqhjgbeda/kJd6IPG7UD7AINGoTzCaG0tWRcs6
clCveEEsgS7Z9o0/HJCsugh3e9ki4DiOc5n9s5+LL5DDs2cObBLGWbPRgEeTxvuRTF3YZCp0QNva
9i1WBpTB2TuhlVMAYae+tgzLyOqMe3oQzuWjKkY09Xj/hDfJHFh8sFPC30GD7m214rrazsoaaJsb
+lcnLnbdVIx/vYXpFz60TWHzEzOFmb5nPs0cFpnFfpXIUVqQ97SJ+hBnDcpyiyravb1Jotjwk8r0
b9UuM20svtCInkCJaR8LVTffZ312v4uxKq79PBAP/GTA1ISxsSzrJ8p4Gf8B0/MUCCyie0JtlbF8
3vxepgKtAQU4efazZ6Karv4Q9W9zicaXsdb8MmMXF1uqWMCiPzOR85x419PjCvob0EEY/XMW6TwM
1nXzlWuSg4zJvQqQgxPzz9Zg0qQLxWmgHZ8opW8HwuMFXfvAe2M4d9WgjIJhxw/WkZdoCR91Dc/Q
bp9ERwVLedQXmwSURUFU3FZ8Fbs7hQTWhUAPsoJqD+YSqP9TeLw0wrAzIcdDqQcs/2MAi2kHDEtZ
XXkG2X0xQEhcaJGe/sP/LjZvGXB2Hnjm/3Ur0Q2n4gR7ZT5bVsvOw2OnGmlU7x5XPZKHjmkOoUGr
W88FbSLKNXJkDDzdVOKIgbBsBQQdC6ZJQqg/OqdPaQHrScIU33unVhAJERvGgkAVrzosOQEInBH8
OQvMMkQjZfB5pHtFNbKQyI93g2bRBEb3N9AgzWhoBxgAGVYIbCbJT99mQqHVw8vjWCOcytbVftvq
vQ/GmBr4KeNA5S8DV+e5MIGVcm/kpMERQWIG3bdV3cc7I17Xe3hHWFaNGfCFJ/NAuQvULJ0GOYAE
1L/YHzeWqfP2Xw53/T/Lb90UR1h8lVea+pMLr0ld43+qxc421sDYaICGLgBnpjtKqVgqqAsUf+xx
UFtBniTxgRlf2JNPcZRvFU5fQmGrn/sariRrG2unujok2DBIrjJKlGOO+Tu213xKAnGNI1u02HIN
fPQ5znWWHK2s8oZEhCBAfgcBCWNDYGS/9UiLlmyAyRErk54ev0FS8pX+22vlOHLIOg2hL9zE0z+E
YeQENsNzkaUh+yuZENo/BoJtvPeHl9aakt8SAMZL3OrU1cQdn/wi3MsvwdwnculCJV2Uj209IFjY
013bzFnAo3kxn/mzCV7cA89mfwP+1dqdpBg+vBL2bV0CrC87A3btQw4+ldz8HheFk+LyQbN8Iu16
WFV58EOyskdCYEzl1jCxtO0AKWfHVHobcyT3v/0hS5wG11JLX/qypQosYRR9l0j81h9GKqGPPeHi
VD+lfjsdS4t+d9BHV+DwNJ7v1ZzYxQCdbhs/27qdy84hX6RxOSDOUBkJP/9s4IT/8zAdKa39S5Na
NUBdfmGTqByxKHa7NFlYVCGXSNPtsOxfAc961ut6SJJ0FK2mZn43Nl0fr+WST7kvNL1By837Ee7n
6k7CvrXN4acjdMjjD+184Mi8VvO7s2xs0Wf62fKTAaQ5v1P2f+l2VpPz8yZ/rVbK6wqMnnSunCRO
7ODUAYqDZCtnUcc5P16rDKdb7G5d4CSVqGcFbEAYWCKJDvrsPRau5uQYJACESXFKhfaFCBgTjLc0
LPbLQeiHNyM/rz9FQ92Abm5atmBD+aFZiTduFthEPMAGSnBjKJ+QxrjEKHqBKdXwcjWDkgRjSwVB
sW9sZrAcLGMT3nbd7t8pXFjTti6byTzdVvlciwHI8YBRoNDvrfEZIj7EMhrZOEtyRHXNFpp/94g5
p43nfGK8CdIYDXvm1hv4lfo8KJgtTcVfZgRPTQFZghH7R03zN8WvjhRdrh+6D7tM2RdpVIn1Xmgj
eSw2kwWnx8f+PNg7omVBOzBoFl+wYtnaYgLcIez8fDB2vKiN8jg7E9be0Ijj90LMqc/HL5zC6YVs
gQrbMhOmVRqXp463wagH7aBkJtg/P7rmWX86dEVdTwDVJftlqrNZCrbKH61UQoxa/NEaLytvJs8L
kAh8dSXGQG20JXonjWYMT3mfKLfnq27pGY97lhuYwymIg8wTU9Kmw0QShgK+e+oBAhP188pLeiA9
XNoRSdshOg1SliordpukLPREVFHKsLRZyu7unB8IAgALT5UDa4/ECNN/6q9OOmorLGYiNinR1IDC
E4gwR8StQ1edpkOxXr2gW+GD1xp7oE10Jsn6L7+gvdSkFrflS8IcX/eya+HktfV67seEQiaTRcYJ
tweUXSyDBi/tY8lFw7iN6wdW2fK5N881ipwzLfbwgH7Kn8hONfb0SsOIW+3aeuXlO7Miyl8Yg7lr
z4UrhB0Ks9NR3VkVUGkEKTlmIewhfvY05BQldfXkysJ+d+BHi3yYV1gz2e9tAcFwWuKM1vInJLBx
ZCyxY/NkwmtDnN5Rw/bPBYSdLvEvSbxODv9hy00tVSwIRRiQ/l5nXOPk2atDo2p6InpsVbcJtMJu
S3+WCO1gKfKb5mLgp0tlN3ap0wUAssYHyV+I8EEPMQF8bYo=
`protect end_protected
