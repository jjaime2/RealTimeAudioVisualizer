-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ko3Klk2lE+/HRenyfeIfbnEB9KEzqJAqp27ocv+kuwJTyJCIpGmqA6icaTFz9jGK4X+rZXfsTdm0
0iFpBFz4GK3SC0/NMwA6i5EwmdcocNLbMWN3JBiDM5+5QcAm6MOKaFXyfs68eWNATTGKBsLjLiaw
P/1VJpRhVmMET/A128Uz9qRO4P0Tz3ZMkqQNE8M5Ub4+sZrVVNpYDI02N9S6lq1bH2w/1DRpDEca
v2e/8tbNdYCmZkrt4QwzaWaWuH7lvWisFXCVV3Zyz/Ftu4zk2y4pcQGlT3Iyg95lvb56IT7HFNI8
MK/0INeVTaydFgGT8jLzHE+Ug4PfBmzfLFIX2g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20736)
`protect data_block
+ZG2RVArUEUfN0aEueJFKU6iLbKyRcxcaVoq1XjL/q2e8gQjrKIf5xHHxp/SbKOFVlerltCaNGBy
V7HvA8f/Z+wtwdIZ34LXpVnejRadu555h8kwc4Yy/rSmZhYYsNMAR//W8QipY/pKIplUEhf60/J2
a5dUtUh1qQzSOp4iat/2BZTQ2Rt0ZKpU/yOtd/gktusxB9dRxzdWQYi4/K8fSu9lRALm5r4NY+4J
bZNVeDRf7+AS9fvpVwPkwjT4ZuoR2QvQE/TGTI+yUTy/znOAdNZt2FQP8RqREaPel/BLa+/JQj0/
J1kz9QZpllgPmUrseXWHUIIGu/JPRvX+FORRi3vLWlU8X3l349jMETlkdkodBBXzrX3y3e6z6lUF
wdwJJxGnQWl4YNPnwo0jVXuZuYF1NWS4WrWpAvwtmM7DFMFBu4svokmgEynkzCBL7EpeS6VHphPd
aD97iQ1pDBTYtzaPi1rqPQEOfDEw7D5m+xKaB3f8w4fXPaQvH5uFjFLb8+1J43Me+qtc0JP3c+Hn
65n/RqA0fEkY4FAsG01v4Ip8Y1Yw+G2B4z0sDXkB4URoKVBmiQzhE80h/lwth3VxZdW14ncvBHrh
p3ilHDDsB7NRGBZ3k9kyIOF7JjrsJIdZMrZtLrwGl0hJKrhupkcZOCbpyujh5kgGaX6mwaW+tcXo
WS0Urt3ce+CmROoAkQQGcY0zvyNGIechog21AOHSm0fvCu0QbuVE/3Iw06KENstKsZm29X4Eaw19
52Bib1aQBCh+bIbb8g5hlU91072uFKxrAdp+97j/CjVDDPatk/o4e+A+TD0PgGnZwvEWN9Bc5Dow
yS6zXh6rR6THt3opaDVxhTvV7iUl1VXvg8bhjAHCXSiZ/7IDTWDmnr4L8VCB+N2aIRp7BD8JZg+B
wGi2KbDb9RRBCeyGYluCCQeT5t4zBW/tkZx8R7X8nGp1z0MAL4oDoYiSON1F62kYUwiFQb7YLlvZ
qyv3IMnBk03076ZuHmQraFyLykOaNVA7br4DmwQ4VXGqu1X88tC12PONnz9dLQFDI+ZreLwagutP
TPcdi4AanG4oBAlomn5tZzwwpT8HR6MKOWnbMcgHYPU3SClcFBP8PeOVrH69Z/mAXKVjy566lNqY
kmL6I4OBhjmu92MgV4JslmP35cty2ZeCQ8QwUvJWK8M4TPXFysiV/lIsGw6vhb9d+LaxwTl9zXCi
kz0SkpI9kZSiy2fcjkzO3XPwPY5q9/i5J7H8CnsKxxQtRoHjqPVUEbnutEK0i4JWjOlhZlTHdpvu
a6S8oW8yX0g2HIll9UsCYPD164ScWO2M9D/QQfbSOr8qirURW2/LIyvxWAt0+XZ/tPjoSBCmmdxX
gE/1AsNoFTPmjWqNqK3XEsvA8Ci3VUTaLUH00Nq+pdwgfQcTAKIJcsSgRzwGC+l9T7Q7yC7iXsgo
oaQovfImX9ufFb3mXcr6OebN+Gau96o/aA74G5xSZixZRw7kBQB3kR26nNAvJEDwea+zfRBGPdUR
q14kL76bWvB5f0jzN6O+NTWUquouYSDQtProMCT1nRSOCfP03hw47fZ1euYL5QmEiq5G79tN+J0G
4qJ9DPjrxu7+SBsf0mFHBtpiNRBw5JaZID4rzgejO8fi1CwAdfAnBiwQ56/PTq5UCellLVTE4Dxj
UJiZrdk5I9R6CoowMXptnOO8suehx4j+9HV/Zhvu4rYnaW3JtfsXvdstsWjrt9lu7u9DihNfeRBL
YVo9A7hL+y3JDoJzfbdiy0HF1ieNi1qB+pH5nQUcA1IJI5pO2oMIARcrtVA1oRu3QBADD//0gaU8
69xomdzg2+ZHMvkS6ubUAZyp6+tPPU0fTMSipluYn0FuhniiUBMmXTPv0p4HCPcrWUeKll0Vvl0N
KOqg5d0Wazt6puFWNADWQdLfPtf0egSiVhBcSePNIXBBLpdFz1FKLPfktI63qapl3+3hTr4bUJ2y
9gO2XMlLCaef/EIzQpMUcPdZMNhTX8A1UhQPkvwSwMuoYFzoCunqxM/XlkMyIr4Od+sqmQePqfOL
o8/FdVzHmDRqH+RCLVcUhODSoEWsOZ1gyKZM9w1WGTSUoB+EwzKSLUSadyRDLtFXV7Pay1YP3lNk
mRdb4onfABJYruysE9cuTguPBsUSKq98uP1jAtejLivsZHGiaAXpczUaGRFweeaLtI/4zP7Winch
iQ7QVh+vxDnq/xhOH8iHNLaw53tDG+ZueoVnVZAAlmPfm12V1anG7OYkoyIf7oCAx7wycGOKoMWy
ItNoiCy0LYgROcCljWcvrp8jnrguh1fssyOlj7GbdRBtxw2NDpB++rVWOXfLpmswGbmQkvpPYHnW
5wDPZ6FT4+tF5VnjJCCNaSVW/1MZ1OmCanQCVyG7lPK2XqSapTJBcSaXtEs09oMcnM3yMUpsQdQk
qAqo1/PtSMLTVldhJYTsY6AqUQstQZr5rn7MldhJwM29MDLDs5NOLRXrmFiyvHrgM4uaaGTELMb/
X5pf+Vq+2LE08nY1eSPi5nJ0LbBUhl9hVBMais8icHqgunUve2RcbLLkshb0K7pFrwQBLZsJ6UHk
ivWLPzOsaQFct8s8KrO9VsSeq2KQ6fTl5XjTF6HmSgVVtS5mJt3tDLWdyrKjjmDKprJWU2IYoPrQ
gNKZv6STtWCOWma/X8SKQZcnpZg4CUF2jw5fMoIVWXChLwoXnDI02UNXEnzpKmolYKt6T4+nnxnB
GaqH475catxGPhuoUKNKRuRXQvqk6WbzgcufhD9TcWtIZlXH4IyzqG/Dbr+b6RvgPISjqi5cxrBF
L1If8vRTsapidecpUNG1wr+FTfdGL+6pbI5RvGtOfntDpsLSGDl4M8KEmMR7wJHG3MY+UaJImtBc
Mc4oszDY8LqsX2we4eb2RABLoFdISuvXDNxaw4CdL7l1CYaKHAs2GK8FJjZyQ8C9XPVKOyM82TFk
L4+nutYOLXfciu68qoGItz6G26x5r7PAHY6hS01Qfe3/YGq61V/1PFoWj39CEv3tBEE/XYzW/uFI
cCVCjm48GO9ShehUs6/8+mYTVSObURyWurOxDSP9ScTKC14YJV5Qfh5+D3FIUqsrq2KpIUsCgViM
y7QfwH9f35HfuaMZKy6LeJZ195C04NMLondRbz5jtRKfZnv7s+gRJxkuhiot61VA8NIxxJZ6PqVl
AxX7uimQDp8VmqdorXsqoWUX3aItzRFUveOgPbqnnxNSQECenQHz27HcRmTKyt8F118OO9wZFOpR
0NYlY+0LXs6IbgcQfYvMWBWFHURJGVY7azoLksq+IO9Kwb1DhavZvEH2LYv+HM39dBt/FVMQv3J4
r/Y3zpQ9gQ1AW/Rhu+m95hoWUPklL5FconNGpOgWars8AmLI3Ji55I+YfbvVfgLC/M0BTDjH7+L0
0Ux66rHiv4CnTJKXX2vxpmSd99I4iYQHucz3GkzazyV6oASq0VwMnItskJfoSnmpolD+qG4XGAgN
sGFyY6voxJybNeGdRjKh9yfxE/QkRWtAcf/PFPUZ6kU4Xo6l9duHiJpv/TIvwRXc7Z2E3Cny1pvg
2CaKHhGeQABXnFsSwN1UbHKbfD8VXjz5DVS/8YWmcOaBwW1QobmzWi3Wdu2tFImdL7Er1842vRBn
1v1jUvM1GGF01Bm9+Q96MKwByFwuPPPtussAH1+wqQ3Khmx93CPAdcoW9rCjeBYxjo+GV+3GdZGe
bfuO0P5c0qozFutR7M0jTIWHh0IOKJK8Tp4cLLXL+w2fJ2h2ccXEp/iexIn2SzxFuLT0nEMyg2VM
znBqqlnVliPfXp5NrGphtevyHDy6PbX5NS6tvujDftixRX2UvDGa8sm1sV0i8pjn2zDVzw4XGfdY
eV/NSCW1tIBxfR05y4QaofAhNjcn85zB/2sDVkbwTrez6Kpkz8+GXK6T6FOMAxDPj4ihj940kIbo
OocQ26o/9Yc7rqCOZkDzWM6dlKHm+82VMktUblBulVhwvcZGaEbNEBjf0WUOp5FPsBIlhNLB/T43
FhtcYi/DGnxTEd8RVkXk36FAT/SoQbH2C3h5BPFHB+u0cuvumnfab+qeHK/5ejoQgzDDzSoCrnyB
SK9dVw2Xfwotn04IUCjWrJKDyDpIq6ZeBLHXe5kZsy4S9aXIz7n5Vwa4obwvZZZOey1rwLkJO/ep
bevgn0XYt5wP5S7dhWxLXV+lxPpE2OnBzlDVliXRFweF5q1xLSuY2N+iUY3NWJTYYWqW8JuTVbun
5759iFZbuAMe1Hf227sbO9moYMIlnRrVH7maLZP6Sb9NDujaJF9jaCBEBUwSUbNkpdISGgPx0At0
364nZnH0DWnc2MpVEq9tzN3a+dIBi9XNP0B1uccar7Oh9156nJRb6Kru7u1vPBcjsLZ0E8f+bZ7n
UpoaTZKtcaWSuOlQLYLEjCkw2UBXH91neZaJh7jgVPlTEE7bts6wiM9hao0oOuGyWfSuCn0kEqIo
oYjxqsUnFkCO/XuUgxn/VuwEiqnmTQUpN9rCsNVDWOlIZcOUgqxBr7UhQgqxA6dtlKt8Kbg1wuld
1HDaCQM9EGGJB4f76W9VbijMRtKTdHkaWPc9/8iZoTr/fp1M0hKB6KExK6SLdgaCkFEh7PRIvX1N
xTbW5OSeCTDlTg1XWAOKKnJVPKaEoRiekPv/7HWYDwV+UitKyNmbpvbfPk67cKWvIUcNlx7jBPFv
VIEv11ApRQOzPO1wwvo4K4XzLl/Xi6Jq3iucsCNbUbKcuZ131adWPApZTnsp8ImZqM7PHRpD3gjf
kbK9/Lddvgsu8A6PaSy18M7TUmEj+8ZNk7ZgD8lVXXH22dSgKuMZW5wKw8s+IPHsQHWOVrDmYS8W
JsTqpLr+qZ9417i5KzF+/WiuxtPicQwMOdPib6w3BsK2JYKpHATtggq0fCbALnrjLMabwcNXDwRg
UnZ6yyg3ZJgSUsTqd4mzZWTdyg24TLlcOvulwzfql6A0rVSHNSZspDPyHEhUYCDAcuItUCKvFKNX
VFvZXeBJ4rSLCpS3IUbBjpaf0tx5WDs1KcKVbQtZhkTWDMw3mvIG3Toi6QXHlApBSmMb6W+qHwai
JMPPs8kMXFMGa7Ju3jdnT+Ycxgk07P8YHOeGa2qDThL+PuyXEnzZ9zg7s2z4+5gv2u/nCseGDUri
B5f+bap+yKxFuGUrb4CGvvW9qIzS91CmWQ2nkSoGRNgnDV0huUXsgC/S2tIdZYkQ2OC2yhDQ33a8
e02K8dZcoSz8g5s//kC0SPrHB9AppRQLNudwlvW3IAjtMu3jS5yTPyq7m/Sdh0DhMhrhhTJnuiia
savjU+fCgSfSyDucBxG+iJ2gWK74rUa3Oy3ovB4Qy+TRUklbxQCm2wgcJffXoB93SZoBKblEIB2C
5qwdzfOzYppdRtr/Zv3oy9LJvh0hS+A/+BcHwpmc+GIi5beKPModxiNCjQyfzQeSwbFCuHWGfIK0
zoWZcQ/pEnWijpqJOq1ARx33vwI0D0KRDXaynWbjPSbFaBOcLxKfiZ1cpDmqn0is6jyKdKEVdvMV
CI+I3C4XtWGf26hUv44tXOMvhbAIqs+0xUlGSZBo02Fc6bPR2zwWSUGDWuXFtUSp+MEyWtirvxGh
DF3UhR8afV/aDQRzj7+NLkB9w+irUVYZJPGmvZkPcw51ZEEqKKOZVRdlmG6Nt1LREkmPkY7jXnrL
U+UCYlwSxlVNn1i7EcDD6ohyKqn7XLP3Lbgt2j2SxRovQtm+mUQD+E0GL5LiCsyQxWEepSr220Y3
mwAmmUKNzglJybdsKcPK49TW7EtrkZ4Js2ZSitotmB/Ek2GhynZchkunW4cPPo3XwN1cifD1iOMo
n68FXvvWBa+YznDpFFTOAQ7vAIBe6xNO/2S2Ag5rcMArO5sLbKlg0Sr8A2vZZmsyLqTOPydnRQ3c
kYKXibUmsvpNvZB32hvBSsQVUDcdjIgBFn43cl9YdGn8VhHVsUf/wzUzwcfM/JQfYShG3oBaH8pv
pFjLAaPBjfgA2s4PDVg82s4f6Q4xZmLIY/cH37t/RfonShaQIftD5B1p5nCWWQhUAeHEzr0BgFpd
7bRN3ipnExKAAyuYoyVglXGxCFYfxd9CB6uRXmof90JvwmkNR1PAJ54Cae512J11lTo3OTzcieKH
OvQD3XwEt9t2J2eFSMv0vKTtq74QdljsGXbHgQMPTBnXsbEzHp/livvRiyzldwpoY/q0GeEOb+4A
m2+ZP15f8Juin5dgK7ncVTmqVym5Y6zdfsrIqEzXIqWEoW0KwXhjn3appGOEhCHRgOwns2tYKsui
aziJ484TUPnjzD/Doo2ooH0DZ0pKL0EL7bsUAqNqfPBwNkPQ2lprNUjpXzynRk+0wPAnGLZHvSzm
CFIfhMGwkC62D2eDLt6DsQV5nHyyFUXnX2oPeqz1QrjMvykhPQ2TS0wTPNn3VUBq4vsBPjDC1tRh
u+c4koFuGPCRvfUVSRx+KjY9kPpwm3/Q0PzoyPyBd5IFWn/hf/R8PldsdsHrqJgLEOLb/kh237sC
jMF8SvQu5D14vJK8GeiJbkls/lqkHWltlFaC2+TiL8HTolIgPS6sdS/7zyZbXG/csqqdQr7AqXAx
eHm9l6QZFMfz1OQD4uafePFnMMZq/NpaRyy9gUe71RoSfW9cPjxOEt6m1og7C8u9TJPIL4JTChEe
M2h+2dIPQAO2AOg9Cba3f4MUUtCe8kLairy3wNn5Va/8XSPnmfQZL7zeN7o1zHlTgLQKog+fVR0E
Bo87xu4u65ZQNV89VYVnV2mIGnoiT7DwfKEVGfHDOhm/XuxNIpUW1WXh5NluldDsS72MMAgot2eC
78Ws1azVAXuKebOKdMss3X+BkV19KGz0H/35/OGyLpOyU8jG9ddBMO1yAV+M3ga9OcoQpqt7nLGb
vJk/MLWapaytw8vHjL3ZsYgBeCcLqrTGQ5nYl0IDXgK773l6K9NoYJ44cFYAL3qD5fapWktv/ygz
9T3J6wvmfYmoLJSSR7auwMg9Tk91NFejuy0CYuyakn8ci4rfvtSB6C/CPhrEiqGdN7omchc4X63S
54SVhsNHgXz1yh6GOEZcNqNCsJQqLAZqkhl9uzkhBSlrwIiSzAsF6v7Blxxd7RSX8rzYSI7IW8AH
FGOR/2wR/lMvFJaqEDoWdrjNleOlhFdqO/msZqgqOCQ2tCVxRKTfKEB2V42Y34kFwSZQpMAM2qal
+XlaMuXj+mg1cd+5Ax6s2nMeLEzyUatnhmKXRkWqMf35csCEtfivK7TYPsft/ebdfh3UZ6rb+W+e
eCnQOqFAqJtUZspKBzNHrdZP2nbCdJeb9cNpIFOQfsm+USirwnUzOxwThBBliSvw4K4FPcHjRAu0
6RjPB7warB4EhZPJWxnqA8E8YOe50316Rl32q5kALVpzfkNg0RyVgNNAGieUcXKPL3iKlJQYyjWK
owZey5ZVPkVyDWDvRi9vQLM/PTeLmlf5jSG3tu3563sakZMznzcX2AM0DAa1J0s1WfCt6so/nrJw
CjXCPnKIFDnJvyniIEHlTBQnhkBtwR08Kwvxs+h1XtcWiOqmiJdOwLBGcsnE0E6HWYSlJiK4cCrq
MKqse/bTo3j3loQ+F8vkhjd1xajbKqzaD1UdDvhZXBafy+eNtk/TgYHr3SQ6rTiVAAKuKdsLYlec
piq//IYwZ6QEvzZWFXfBZriApQ8auit+ADsk+dqzpUo6kVyiSYVtUhGy3CE4dl7q8+ve/DaYDpbP
+BjJslDAr3obmxktGUCvUu0fzb1+JN3Z4ACWmBefN0/5M8aN3P2hsWGseWnkqOrv547y1B1011TH
JdxCgmbHbsbIxarO4z0TqWwHgGWwQmkVNCRFlYQdTzU+yG9AM3EiZcq/3Cl7gdAhfBdgSK5QLcXe
03zrfs67AbuEBJzP9QrvVi3rAzEJD6Fr3H/ImoAoov/4ru99IHO94tHiN7Bt2dRQH7Rzdt2ZfgKr
fS/2dVXz0MXHhbkSmCXMqokKh2JpiF52v1XSRVPPNfoFF3sJA41SCJ70inqLi2Pp3tLS7mjQ8eMD
n73vZNEoHl0GsWlxSpaiaooPsMEKnJDmoSC8KvP7HT6jwdexWPJOFhiQlYow/CNWAgolET57DzZr
FDvu9CoiwU4LsgJSQlmXrbScX5GefT8Idp13ufJjIyPouYQKL4zUW4tUBu1g75fM5xGWFBY0ZyXj
wkBn1F/DlFXs08Xzep8zlIcOPFCc2XujouEg8aJsezO2bpJaeO+IGmqfJSHMrM6+o1NhCWUD4vUD
08GH1PBlCT5JWfz4ibX1beWsp8nt0HRY/YWNv0m7wQzwSI7CbIwZgr+SoHyhlBDdV/PKgIzuQlOF
oAipcvxLlZCRgYRnoXVrCwj4Y6w8ZlamKAdmXs05SRadgy1I6rRZwSsntD9HI4K2OUVpkmzaK+7A
IWg+DlsFe13GR7s1PmPggn86YLiXCwY+GQzA4irgwVP1G3Nevf1rX8vj98h6QWzDv+vcJY2uWWA3
SY4zUEMf3keHYLdgRsPFPbeNyqPm0sspMRbzd3nyGMTzbVIE9E2UzjsRSe4mkzNNvHnqS3w8OGxw
UWwKYiYP8MGT1+M6Z0IISbnaOEXCtvwZ7AfsCQnWlW7Ea/XN3m3eEdNA+GHpfoqHT6poZ0i/k+9M
98bp8lkjVf/3r5Oi51pOF0YAKeWAIA6Tz/exzeF4ABbRWrinRDTC5LOgriuJJCR17eaClqvI7sq0
+DEQISoNPvkxcOMsAa3Ueay5xRakmHbaK3ug7wWbSXZ+UYvbO8sfd2fe0e8ItUe5JQPmIdgQFgdP
U8HWuzDtpwoKDYFCKv95gcHze9zr7j1sGxvrFhIJU/JkMO7vno2ud4I2IJrTibQ6NpKa8uIrJBkB
zwk+8FuKvbpUk+0cshr4+O3w1MEZXsvZ6xyDmistcv0Tzy2MH95kAofqyXqS2QGAjCB+Ep3w7ked
amqv3lOjuESSuJ1tZX8sP0rHhC9KBFEeCmynDKWrMufX2F2rtf5KBYF2MbUFZDFN6tdji9ugVeVm
AoKtHVsd0ElcoCc6mTbQ04TVY+Y4u0kf6fn47CCIch3s1rLhyi5W3ruBiu9Sqf3gQepUhJzufVYr
ODcQqNYpYJf7b7BkVt6YbHhGfjp2NIZZIB2eP38Khntz39VOaLi85VljUWzhf427IviZG8y5XZv+
tC8+no9w0zwMPpM+PIyFJAdC3J4iG2Fh3wQk7K7e2R3LIKFjkV3WK8yQAp7rw9VpwhbGzd9e663w
WJFTrlK6MInWwOwaYQjpoXx7vPSFAIGDmjXGhgFLt7iHoLY56PTOfqbCHRrtT5tztsiAqhSvWUlH
nr4b04o2nxm0NDJ9wA4p680pIO0eBKlkStROTvTk7F1eEzEBiuFfQ2jrLZcd39runHsM+L7IUedD
6bz17WJAzTvKUtyVaptn3i24rG+mi5I/gbd//wsEA0uE3Qwun3S24XWpj7Q/6GypYl5lyEei38Bz
4lbTU1XPTqBWGghI4jSkvLj6dudcs51tZ6XLESDdpYfM8YvbNcsc112rDmjEL7rxwSY9aQIvJ8j1
WjevC5iM+Kz8OHBExZZoEWk+s+n4FYzieswBQEGTamftCuMtZx9Oc/9+gHVUx3zjWsDM7MWSoPzB
iEzzJvNwSH07Y29RpnkQLLN5t+z8IOplMS1UfeDPaj5gg7mKXYSDOUC9rCSbq5V3i0K08Ei2UbQX
DAwYcP3obWzWrk6TYuwjW5afoThm5HubpwQjGxkbnBHCX8hnpxUK1RiG/KG/chPtbUtV+hnZab2W
H1TUsWhqVvnjNmknUUFuZA+/EiesKi6HZ13wVvhXh1p1aCBAPV9X+2Q6aPIi01PQMtZt7NV16H5u
cwLf5/Z9aQeOdRHBydZfkgq6+pNG2h9QQrQG+sgH1GH4sFDncswWlyJy6asfqNP8FGCjGg+LVfmn
0dhgrNFpoS6PiPYAQxoL+8Hx/HsZvKGiBTVylHBRjdOozw8B1nUbVexevxwYf4jY0B/gZ8Z8CdPk
c5+fYa0QA6ejt/nJBYiS5+OxJz6Oxoh1OMzizz9eiC2YmMAd46qao9R3TdfXT+BkrXwfsT/BCVy9
OsQBfLu7L6zG+gqMfJZ58R3Y8xnI0Po7WsSi2QnSMKRj4vY5VSap+rY4KzPFR85HpcDd371W6zWi
ngZMszuujoNIjkCvTeTvoZLdJkhQPcYIBOejyclTAoPltdNINQ1Izwaj7v1kE5x4l11rS1BldBEq
ZD8QXGow4Tte33QZBPognjJE1Ia5eYW+tZbXXdrd+wufwz4WJQVel9YN3FroV3MWlZMfUsvnccMT
37YsAMc5ntEE6w63OrJkpscXqgtvwFsf+VDCi+ce/LQHGmEQb85djWlgChmqdWDfDKs13hRb/Q7e
RHA0TYEgZ+2Ymv4yuwH9dDL9s5w947T4fCvTH7nOG3ZiJvZwAUb+/3qLxJRW3VBFxy71LDk3abxH
o95nZh9bjc1W5IdNyDIY5g6ZO5OUeuXh2rMNL4LVQ/UBVZmCL7+MBzbGdgbRfAyGjCRCZ0VcXkGr
7kL3bYfIjFMINsFUdO1cGbbdzUDezluKn5UZKS0F0frS1HP+dbjko9JIDOMMVJHsMZpk5tYNquUP
bxkxuZVUYOFkSEXJMmpuQCS5+5M02UTy62WkI20s1IZkSFxI8Ga0CZzonYoHLZCcfCo8r7x0WHq+
ZiHTS5sGJ/pmPp2YgjMflrrDAv1gvvfcKZ4LMwEDE/A/9eOBtVKUYzr10qkQGud89VCO4IzrBLme
pf69NFGr0HxnIdVOhTYjCdozkLrciT3WMh7Jxj4Q7HtHMmJ1UfY1xrqLxaWfHMXFXKBYyn0UaLCH
nZgOzs6n0lDxlTneQp08M2XwPTO9Z+fPrrflxS6X8tiedtHY5t1xMKsgb+T5Okd0Z8pYxtLjcuRP
ehCibz0+eaRDwnUmAah10n35NFyodKEU4dXTKTcMr6WkbRlaMdQ2wuqEXXFu70tyS1SMd/KIminJ
L4IEE0tqxmG8/PLazSUeLz+0B7wepHelT3/yWgmRAxZNczTFkZBZzgyO/nwcjyDp6GVphdtKZS/W
jIQBVaaz22z83/O37SVGcXZy7ldsNpgrwSyKfABGidjBD9IzuQol5KL9LkcAn28PdpsUPy37OkyQ
wPu+5Hv1lmIY7XU6RbXEBxZus5kTfxS1HTJWbLoN9h5hAwaBgal2XX62QBQpEr9QVR5XX7TiHww7
HHl0HI+FSr6XC7KbmhSSKVt42fycgx54s0PIsuTuVd5vwj5j8MQ22ZsmZU7rcit3ntOM1OGiW4k2
mpB8oOE780yb3fPMSWykDeZzp2360Z5bWhOETHKPeaf9OtG75s7TVLchJ2jvl2YF5HqVu22LNMJt
k9gmyLOhF+30rzw4OoL4nzRVfmZOVJ4XiG9bulk6qjFeriFAnVYlNlR5iV7uSjOoqDWYNZpjunvb
WFSVupikW3g0gKEdK7og6Iyl8tXB3L2D9MQTImhKJsVkeuR79FIr/P9/YU9RInx+C0Fz9GCJcClA
zINLsdDAC88iNdl+rCoh8FRiReA/9eB/Nz+790+KfvUwA/oGUTsjGBoV/ni4mD+LowCM+Y3bd2Hd
0mqEtRkhufChcSA7LzEYasR1sJAWtOu9ayBknS3AuBgURTYcjuBMSrKSk5wm9aC6Gz8kERAar8Qb
YnHjFW6QSIWgPFE64xZqEOqY03AScsHxyMUrXm/MqV7Vsl6Vkguptpdxuc9grJfk6tIzpVTs6A4C
SBp7Gm/omNeHI4um+X1r6SLgPRkNZFODTg5kghxMqkfUol3c9zp6/DiK9fP9TA0Ev/mecTCVpMWZ
/jtajRgFfdfVb3zN/Pcm3V794eiURYMHIwhrQp+g1ejJ5GbvUfOAlczWVe9de4UPI6ikA82cMDXt
W2SOxqapQKYToAixk4jDprybnV/rLTCnZcPjM1X9jhMcRREy+HNTDaqfo3zFT/blA/5BC6wDUKRb
EIJ61kd7meZBMRMxF/EjzQd8bHbdNCPmDQlAjuqvD0NoyGfnbH0zlCXfoMpZlcNjSLDwq+R+5qrd
Mjbt2Zk57xIdm3Bvq1VTyIPA/Zl1ZIPi0RBsR1LNYuxOcgEqGROuoEYLWa/7AecxOW+HqcLYT0SM
sfSyFmVak34cYpBprAOygcn7aRMe4Zii51CjzvuSZrfO/TMzTy7dgoFsmRm7Ul0dkYkBlvs2IzsE
/5+Z9yV/QeXjfncizQKb4WcIcz3zbs7RyjjZOFs0zn3qwETaQHdscD1iZada6GziBRLhDfDFhu4G
VOj1B9nUfTZX3I2zZ615bSwDR3Not5vl4rmCHNiJ9xNUFrOnLDkzDIch/TKcLx/+w5qfnDWToJGD
NhvBLhx5SUiKInomLeyYo3xSMlYTVVNkArVJvcZUn/cx25EbSxhHlSIWxGjiMDkvg+ryIA2hgRsp
fU6+mABNMcJyC3fxc8/0M9jJw/iGGYWr1OvrNSmg5HwgDAB2UwI9ALe6VtoR93n6WgGgg4Z1cLzI
hCeuOnT8DGv2rn01d5uc1VGHqSzoInE3lgf7QLaHICnDiCWKSzcVEw6xnavGamJP5f3fruKMDEdK
hIwOrchGnt1oYax654CF0w7oerpguBdpnhYjE1NezP48tdJ/bWsmy4yeDsYI0MBcXtamCOlZOydH
uIW/icFKrYHGUzaQT6Qsfrl7iDvRFNJqXliMTelWVr70wKCaR72iCULOMWerhoSNBFlelhz2ZXTY
TYXRCiFQOGlzXJkip7Zvm1qWveX/EsSMzy28FveK168KKoXrsE+r5tfc0VsDrEb3h0n/iE6d0Q+v
HDw56FeHT79tItcUWjSmTxp8v3F0tIPm/1wjNhxmxxx5UDtgYYrbCxv+v2YBnAwwRIoHdkUr/kHw
yR5v4IT3eJHpY0mdngkfucKHToMoymbCt/yOs+tp/Mx+zE/pCW7MIj7aQRH4700pO5HxhPjRnF3I
2P4I1ZwiVBmwdEugNshIa+Ypuxh371PoINxCHjWEmuWdKBRIRDYfz7GspwqZlbE5GxHGZhnycLNk
oQUVQtmsPNajnShlGZS6VToLjYMNnt1a9rf488NRoLQt/XpsCQ6DnaL8cuSUUh0pZ58iPo0EIRqD
qGFDVGkP6tflVBbODw7eKbrzTrBNxxz86uW3YSjLn4qP1Whk0qqlQfmrXgN0QSPzdeR8XBUbp1hB
ATzv2NEfcACJBrWw8F2XfWLFRw3g6F7bnZxL70KagVF5Y3srRAdcZgPCi3cxmjzBqvNZS3pCRd6b
DFiK3yJZPmo6WQ9FUhsUsqwzajboqmXL13r0E0/7qMZ4qoqHukl87O+JBJqlzODlBeEy65lcQmlu
bQn5eEgsfw4wG7OwaKxxRMD+So2M929ZHOhRj6XdHT4hJPmZzuqnD3YiAdM/lV0+Ww00PblQ02Uq
ofmclLRtgjM6tokLqPfLGdKQc/qHNeAexp8s8iB/ct6ZwSmVTuKQveRuoLpyzICITg6T9VwgjE3Z
ub6sQ9w33tPKFW4r10nW9KYsJcAJXQAFpk4FUsemgsQDGIetSdLfmgZPIdcG2ZZB6z4Ws+v2ymVW
Oc4b0sG9Hwt2INybtlyg8im/IH0BD3ATH6AZ6l6cbkoeK47sprlAQAh6/U0pgnTygXHphwq9U+kF
YY4eCVtJsoyz4wjUUdGd5I9dVkApvMHax4ybBhxeFPw2qR0AEsyzX1Md/M7KSN1OVIN7g6elhfri
vRFYklh3kBp126Q6N7aheWhCuTi0U/slOJ9UvptLh05p4xv9seBki8xqgp/F8O4OZnBNKCPiX7DD
pNU52qUsus20QkAtf1+bmbzgj67g65mamUlTDcM7/0oMLPkWyAzQzDEt3sETixxdMMmGUj391OAv
5iD0VO+a/Rh5hUWS2+tzZ9ZX/U4qrywZE9MVc4V/dxTccgTcwhNBLySOMBA6lwKImqKZj+9qAOJy
LNOV3KdMAea4iBiqjGkwtxishNb3ywYyu9XDEH5X9ZTNGU5eV7X2vA1oITYI9Fp5xAxo/FOqop1y
cPrjhoqjfXmZLpbQyahs/8HkuoU0vmTSPaplBFwzxfc+bzY6F78yGIVyRSReOA1xFjMXtuB25M5u
B/gRwY4krbPuRpx0UVt8nPdRl65RZ+QAAsRDWgGVluuR4sTJy9Z2NqywnaKcK+TazF++HPka0sCV
bEJ0Rr4VCma7+3M4b4s8ly5oH1SgC05piHZvKHG0KOg8sUxdGKFtXLcmBkx8ZUNIqCM2TTMSGmBT
vuDPTn7On3i3Ajm1KuvqdarRN8s6bO/b3bBOcy77yYWWGY5hRVxBMVy/tVWgC2K4bgP5OHpg5cjL
7MPTm+cFppFbG6de2ugkr4tAP3UBHC1Ym6+swC7J+xwhL1vj2/HEObtqAxSjRpcWPuOwmImhWwPm
EyrGFDhvA3gFK5IyqF+mqeDCkKuqPiKbbsV8WaOJOhTBof4E39UT0ZRUjYaMjsMj6iiM45GmqWD8
ULPYUErdDPYUAc4SG/CbRKb0xc5g+il5DAaOityL3ibECM5GfgM01PzI5YDgGIbA3++GfYJdBpD/
47vl92kFJ8qbr68EC1ae9UbXkUUfYKuZPUscsEon4CZWJxhsgq24i6IA9dQWClpFSaAKOa8k7Sx8
RjMha0+7aEkE3IfBk+y7GQWAyhJYQsV3c01Ze6qxcPmyKTMYFV6Maq53PxhKVRhk9lf8ENTCTdaC
qkZkyrTcAWCMl14stm/eOVHJ6Cv7lM3HvNEYAfCDYQLs+cPJ6VgnnUnjFqbbdbajOofvtA8p8TO4
QKoEH2W96A1RdeXoKfE/fIwFqoQ7VAvOPrwABSbP53NrSXs0BISNWlzea1jFud4iiINFdAGEc0x9
Ga5+ctGB8N0tJjScVzRmSrBdXD9Vu5JmIG7Mm5gyQcSgIyltOkIjFRpeAXTVSOIyqPhN1PaEjVhF
PpRpJsotVamlc0E6MV9mcqayxINOOna7u0TRjROj+MymQ8hD5CujI99WnVuTa82s/mBKxRMHx23d
tSgVN2xlz3y27su461QrqBeNJ/pgNHPIUuCZ3gYR/cdB8RpEJ7EH+Hmj1+GtG0XsD1mt8q/+w7b+
AaPiokC0cnvvCHZZuafZv1lqUH8miNQuaZ6av1OD3/o1mrS+HeEZkUC0LMeDNcgRqMmVfsncx3VS
+dxneFn5o7xe7Da1TGu95t6GnEB9Ac8AMwF35EHS3FWnpBUkr8Xi2WpSDIPLFSpxWk53IcS/0HNY
LG9ffiJmQIlyWfZSxRfcNw6fvILbEeNyMuQ/OlYdlbuBrcfYH8jKL7+aHWJRLrPqRib2Ptcql2W0
DOYpf08YKtljwdjapMi8j1tUe/xYsDIgWhCCiu0idWC9GulBmHdUgAPPAkJIy8kvsEUur9hRbaj4
5CrUWSbngWcDKbH9enb9Dx4GsdcyxuCff0JgouQyASY99wz8/rz/PB8k0L/qua1IxFUjt3BZo2xl
s6q1F9q2/YxftEcwCx4TXuEhN09vroVtEW8yCDAupgQhIUUzcN/ARF1+NWIMdFUoYa/GbVGSSYbE
KNnWUJc+hxyWfV6J7ookdp3KJeNAgmJb66udFXlHa6yrdNXh+vJUxYtoNZoka610FNQZGwoVwXVv
tUxWfCsEb71dZ7/0fZ/wOsd7cCVVTzu3Ch50oOvAPS9DTWLEtbuDS6rTwF0gAfD5UMfClSli5FWM
6WoxW2+ufbk8//7N1uP/3nB+lrTPBovQ0jHenCBzlj1oJBMzzvu3H5/LoSuT7eSI6BZ8pmUX/hyB
p0a0HsAHbI7NFxy3pUY5IWEoKtvsZbtzXIShyxSYzXvJ88sZuf/9ZIuBgxXXVKle5xlc5ykHqxIo
yBW//FPPA8LceeWVQ+XQWMDH+utzfCSWtuxKbrzuM+SAPxs90dXAvo2F0CyBznV6xi+s4uHHfxiE
zwKNnn7cX6yFbHTcl0CSroVFIbmoyMKoy1Lf1sLz2QdG73QRXHHyyp+/w/V8UTUQQYtbAZELpLKa
/iOqlV4FK8wOcTwDSWVdoFsscF+ocPIaRcWbTlOcOkCULdA00GeoL1Vr69GVX2Gxi7dWqS9rGALa
3jyXMibyK3nQbqDwmNsaqgmSVpVC0rwaAzC0g0V75van+U+8vshNLRXXDLT7/jj8VoBKzOFbmHh7
w10TKCe9FwsO/W55rnoQqayOOUd9N0jKBmZmMf7ooiKpp7+T2+W04jAUfM0zuTZecKokhyclVL7J
GOdmmE1Aci756s6HmKyuX05qTnjyzK3TfwsU03uaEpox0T24cSRbBWG3nNBpwuJny8PatX8adaK0
995Pb79k8knRj/3heY7y3lKT1lpsR2u15Qa9RZtpncQYCtSkKUhN15l8jUqQzvZ0KkINUE3IOOe2
A2G7VSTjlypwP5e5pu47qEIWb2A0aP4eO2hPMCPSuGBM2j1KgIGwq0cK182E8+oC+myz88WJO1+j
B9QfiMuHd5r4hkaBG2TFr1MMpLnHbrbF1pBWNKg3P3nesiCONrE287sDhVd0M8S7X8TitQcU3QTC
kFjcoFpmPgnaaShn2z4SIVaAe6x3xFzYsZhCuwpujgeB962OoYfYmshraFHLgRSdGZP8GTn+g5fk
VoN8EyVAbVu0I7XaiRe7ftgJHZIas0l9+VCuRJi8oWSZzRG8hx8J7U04hZfAp3D97X0D5age/0As
bWJDIzkgl5nMF60FHRQRCZamddl4Lb0d89zFSDnqQbSkk+XobdZXt+TD+LEyCEYEYlPlzJozx51B
DQ7FS67nsHO8X+z+c06KOXhWvye6qF/lmWp2RGMEJMOte7OObRYww3Np18TaSKxdXlR5Y+tq+Yjg
QDCon/a4MGsZFWBm3ROFXwdtvtHQL22xLXYNZWbZRa5qpi4blLlcZEJnRPNaGcgwtMMU/gRyO6kc
eg0nQmB8zvCK3OPsTRIAq21K7GdB99oJYJ8CBTf8VlCR8oX59Zfg5UUL28xaE/OrlKES+playMi3
SHwN0cezhZqSBpUocyNZGCzEYZ4ImMhqa00UfkFmT8kgftsqrnFpRYvql0rYamY9bKPLVQ0FVBLr
iKxQJhSNJhicf9WkJ/xHOpDqAJwi3dOAIMBGSimBhtSWiuNsDbIo9zWsMpCg18hzI7V+sv8+8lkj
2Be4gubWny5DxhYuhqeMss3mrhOqRR3uZ514tXHb63c3MWxcX7Dmqu/tdA77F9l3avpud814/sTA
XDMQUpUpHZWiVbjeMiR/qGvd7//zMEXKqK+nVGjBxzREY1we2AldE101eXQdmGCtzvshxiRHYrWQ
gKqV3stI/uWQPiTrazfJ8xrJ9M/lyhdWNE+WFUMceKDpcSuLNlLxxJ6anvwfDSkh3hn3Ne0WneLu
WM/Ru3kskWF7yJoibHXL/zvrO2pCIVMICuVXxm0z/H7yWGyYBBTa0odTgsL9H0m6l1QDW+OWSEMa
5rXfCx4FKZtdrvfoEwwVov9COBoljhuhYdsfOWUEYBBgx7p8TLjcAtevm9t/MDsqosQC0R3oMBUG
vYFPjx11xHgMd/Sr7p8ZfO43ERNsh7mUl4aFevIepwNRE91p5b+Gx0lDf8dT10huTFsoco95dgbY
K3+ziRV2/sy3S7pxzcpQdsdZh1AezQf+z6w8WXUOXZ+MFAqifXRgyXNmHLPn3VRgkUMKfpH1Maee
kMrWM11HHl4rCEq83FnY6Ky0xzgcVUt5ZSdRUw2wuIgm0bpUQWIZ1US9qMfFeA5o4hmvC/XSxgu4
K0Msz42+B1fJcghcrSh6MikQ9v14rWUDUHe3Uq+MeShHlc0XxuZV/JUdWecVTYEtxf5DJaIhPFcG
cLW+hGg3o9VFlXjBnYGw9M39TX9oc5AuScBYRnxoYlkooCVbpDQUOACGwOwA33QVXXXEW+ImihtN
yVcguHQo1xbWqI7bugT/WbBnU1zEew1yLkIJbjNH6Lt52Ge2PXlb0ONMYIhIIRIfpjQsCn5UCASz
9+AnZV8alvdb53MKiyhebbYvpnmPfgR7cenI3XDi9JxiUnz3O110BYHPrpIgyLj2TjOu/VSROcjD
MGwRiEWhWD5Zl3TS+dMNMo+FMAsD8DlD0i9ckfevUPxLDSoOaPmxILSm+2APu3NzTB5Ml+S0T+pH
Qbtc8p3cdv0kLD6QATSiwZK41yPiEWaZ6hbxJChHS4wLlwOUMroShN60+fnzmPRe/bMzNPjosiDg
cb717+IM0CdcXu3dpzzVp7kJnHStcjqxl3hq1wM/qo7ShB0+Xyt8tn0WfBQGCLe1rVT5U+mFWc6/
4cC8Rh8IaZ4u528I+xdRHZFVd3wvGvQHRKP/Iq4BgpkvgZP7LEv3B4QucSIvfwSCELW35O1fII2h
iqIb3g0FCTbT0p8LtI8aTrxzFH/l7zXyceBfEBN0HjSTihKSySfuRHYadGPxIQe1X77toBrJFtTp
5p9TyVrXS91GfDrr2yqsaV9fxME14mNCz31dP3REsFTDl6I39xBKxjRrh2oBSGqeyXNDQaLkbkhe
46StndQtOyS0JHBU96xQkUBBzTzSPvUzEy95ksgNiYS9MJMRaMPIRNikSRf27ZRFrikGOD5ujM0C
Om07KPQrif0h5Pm5BJBG0MIYO9pCx/q4hkIieLW3irTcxUmA4vZnX78jW1pwyLFbcm5G820z/cYt
l2rW/efgWw49+lmkyg0GqFsrka/W/fYrhhaXaDm2F5sbCVSd/9UyUxXmtMWWdxci6Kh+5HSK/qD8
tsosPyIRfBnRN44rlyw98rK/vpnAMVsB88PCIxH8/sDrlEcB/HMKJs1Ehxqf1sGaL313XcDETBuU
cuznm3Od/vaHBDSVW+snzoX5tZo9WlBFZrOXNn6kA2JpM/agnoNMiZxoG+d0gFqGiznnjTVtkzsD
K3TMgSXWC+UVqrH0wlc+WuPKl0CzipUOomoEw6/pBe7KD4n4My9SJ+bgVpwWAZ2XZj9UmtD57O8a
16sQNAMgRYCQeIk4/jN0kUTJCrsOovOz3C/Cuvt/qfiWZgthuBgRg+qwPhw9E5AMnyaqLs9vY4+l
EpjUCMQhSs1Tnap9mq/op3t1EaqRRLxzsx4o0fDkKLyuei1nlM0jUzeUX5zYxK3BXw3ZT1RiVI/f
qCDuxgi5f2YVyRVK4OzTZapnxorXfjXOmQAkDwnAQbO9GYX4fRjxs+MUu69VeuCNw6/Rt5QY84kD
OYc4rY22fW8tzJSVMGbs7nl4iLB7uEzpewsX/0DUY2hXsHc9605sW3nDOyrANRLOmZp+Hj/Fd6Dp
LcM1DXGdxIhzd3czWchowFbyz0U5n6YCQkOdL7JC51K+mjQ8JNlxeiM3pjFA65YGrvp09uSdOXwQ
nWPo7nyT5HqNSEd5/oKx9W62tt/gSGg2nXlF+yI7D5NL5QpYp4B0fBMqF09u685K0dflgMvs9Li8
3swpSNYfxIItRTZCUY55IM0GZV0J54tGods9R+NnM5RF5IsnAlXneAjaD7gE0LhjN1ezT7XYs/8P
hkPqFvEvzkJBKDy1ZiLY+xIaYdUh+3IDORKCpPtA+3IxZ6e8vXJ+I+DKjX8COfwjQQ7TWox8TEhm
zAonTY86AvkTTSw7OgHFnsuk3wGss8sDv9HRAt55aq9CsRuf3X5N9WROfXfW2yvG2YV6vmA2m/AZ
iIkjRQltStAV1727YnK8W+fPqcYqxVwJoSmpc4Xb5gN6xVGssTNX5Ve0neC10aBwiUnZs8txuqtO
vtmIEEx7VzgNEOANf+ZwMDN+aMPHe//AvBpTneNP/G2lJML0RHGkPd03rH8aiSKC9MdOfSVBJISv
9P8xPxf7lSDCZPFYXJ0MPCf3SQTy4cj0Q5jjf13e25BKcqH+BS8OchVB/1OM1yUuPFe3kndqoncG
7ljDCZL0u4ZV86cl/H4XNYxSNVTSGUYaWHnUqMt4xQxMUpMvP+1CbXXjR86LHbCOSxjJFx7niviK
gfnu46gBLDU6XPl3zvavlvHIimEzh8GkZnhulEDEaoW/tB8YG6jY4LE51bI6Z6WbJDC8fnv0YOd9
WCd1nYmDUYAakJOeTuckyo16pjxQkbbUULKariUedbKVapFLR8aYBEBjoFs72Ii2EZztny6H4NQr
LINHEnFMJtNgho+48TalyV/tRjxZ3ENkzyyATQ+YAJcNL63bMNX43Tksm80XpK6uRZC+oUzc74QM
MUzuEvHBmZyh+Ybj4AG8eNO5ZY2r8uUqjwPGr2KE3Lppl3O4MySNngFtZX/YNXT4y0IW4GzD2SXm
6y1w2cRIPhT4J7dvgoe5omh6fXh84udrypb7/o0uz2zdYTT/wR5AlyzQ/e+LFmvnkJGWu7o0DbEE
88xoadcoUAIsLfMmJ0t980WccrxUNAvtaha9J01Q3CLT1o9QtYQUpsl4aPGrGeJFsumiw9pJTfWH
8hTUAapQVDe7QAkpQcSizxXO0YV2zyo45QBYtQwkMoyNvezQyeT7sEr66PZEGcyfGpFhc2uBvRne
e4umimQtDDA/HsU20MhCDa/tAXp6lHuT40sv2bmqa+02dIbQgUWW3GnsrYsX2ld2MwQmOZOTQwq3
b1k7d7gng8HwSNe3AlBb3Ac1yoo9STT6fgPUj2etvNSlEsZpChA2W1fXPJ8uyIwYpV09d+LFxPsy
5w11BWsUHz2YjlHWRW2SBqdj6UzWj0/LFsCa/F04uN+dAv4b8YSimNTrqsdgXQ8HP9GrSiQ6qbQQ
ZYyzXVo9ZCj3W2DxwkkF001B9Ksa7IreiheH1EA3ID2SroBJeFKIGc5ORZWak+yJTZAdwXhaVVYB
d6jPORUGzlgzt+ilodzl/SqbqvIY8vVcC6jpR2cPtIZrsn1ZI4QA4p5UPIzAid1K81rwjtYtYJow
kmxUXL/GlKbHCaNHnyYUC6pIskzYIDYw9TYTIY2mvrKtUiTTPP924AgL3PNWTRERbNi+jHD9cRZD
PWjKW96hOg9vgnBLKFjdsjoqacCjS3pqf/eJXTypeY4mb3dZgFNEXWobCw88ho+N2YIRQ49PzwBc
KK4Sk5zL4Tpcf1QbR+rJXIkfVLlNlpynFQgi8jRx4zPvx3S4GW0vHJUphoGa+w8tmr2wxuKQMoM4
lVASOG9Weokr5xF5pb6Ze4AArVWDdjfcng6ZVZVYOxikP6uytWtPV8e53h0rChPeuXt+7unfkJpu
dRLLYytqsnr2cDuOFdaMCCMqd7Cvm4yjDH2COQ+pGsuwt5IPPHnmku8yZKSONabLhMk/OtUTohJ+
2TmroP6f6RzJQKcqyfYiv+baEtFHdyZ9/SG3+DFJCBRg4lGfTGW/er3gpE0wpYq2XlbZn13e4JBL
CdlDjfi54gAYw+ciJgWh1/y0mLFDHeHFQ3m6LyKBCQNiI1cmxNF2T5T+rcUBBcTQ+Rq41S3nPT78
9hhNqPWiOzRaL8uNnDSbW0j2E8bU93YyfqgxI2q1+UPWRH87sIDUY0OXbDJYZ01npH27B2XPzhTv
FaVGircv7D+vHqz1a0itPXAkg99+DM8Vpg+qtp3V5CRZjG2vlG56Tpsjd9YBwaYhJmH0ZfQ6CZIR
JgbVP3GoH9mKPfoIohEaBB/xjMiZ3OdJ3JM18el8mONZrkNtfGF5mB36EY2Fcx7qX2t2KSkdLP0S
iDgFuQiZ7kkGebr8FM2q/yMs2KUJ8300Fxi4o8P/6bzEzA65ka64UTj/Lks4oKN8t4m03CR4Ycs9
GMl8BfgNQd92twIp7obzmDPDbE/etGbU3Fvc+gaj9hJjzRq7VdiSxG81klSnPHx3DGD2IBHD4QhE
txXetBCBM2EXrZcTFhPM+AzzDxSQoZSRu56zjHTrey8rdIepJN6oEK7uJmWU3FQS1/tvLTOjneZt
HZjZtleL/f/8jooDCfkbkGiiLTkYTGcthql7oBGPuOMlcg+71cYDFYbFftHNAwQsCdzMAC3aecyL
ehzBs0+gDgxUGGiYtTuWPJAuIJGavlTo4YnGYvLOSFzWRcbxdVhD7C57oZ0FpnfjITYoHQ3zfnZs
1/j0FIX7hr0r8StxHjg1Hl50RQeQgjh7ostSjL6BjJZMVaAIIeaEt1ORNt/du0r5SE23MjeDcZke
hACK1OWJoyciGpzwdzI5aslu57jqxATUsEHCcY1nFyDKB3TL0ka6Nh7xLXuDuOTYCdnHrFj9Jv0J
LWGY6qnPfjl49xnPxma40OSjE+b1ccdkzinOcR4I44ur9D4tvI8CQvaErGgEcd+lGjhvk+EPrM8i
T3NS21pE1AqnYEnl2o3YcF3orn+JGYp/Rgl5u4sPZgpd9I4FbAuN2/6nwgP5HB2ZZ+EQEQd0LIsE
tK3ZCh+x60VNaX+ZKMa4qfpIqvlZ/LZ84WSZcerJWhmh+IWoI65c14Xp7nqO83++pVIDca0ApQYN
8lhdeXGgwYrN4S6Jj/3eNBeil/Wv9jX6MtBnqHj2bSnT7tpmNSFGPE1zYKAOmC1RMhiAQcfJt+7g
mY5YSOoxf7LwkdifBLqPGWEOs378HTZ1NHmgi4cc01CAho7n6e5HZ5AXmvWpgJUzIuhMLr+eix5I
wEzFj/Tu1ebipwVmjJhSEoA4EBWSq0u1/xpYhXC+exBP3Mm9A7Q5rQMmcjbhuws2+YFY6/l0g4TD
Pk1AzwB6S0n+QS/JoaSBgOAVkLvmexeVeoN25s5h9ynNX8WWrWhbeItyi2gC9eCuAHNklNkIkfy1
+i1ztbwyXyB/5XLdz0ESBptWwtL0ViBRnlMvw0NZ2zQMZXe2bslu40bUY9LCCJ1pj2E3ox7mugm7
CrYNwfCviApqE5LMpUp7WN0ykDExm7TYBQC0cu1YisP4UanFRt6uE8DH9slecrSNcaHAAWXIIfGR
UVFLPXWK++B5sWeudnC2uTMuYXL20SBPEF6WGf61f7BspzSaOS2A3kSTqVQdClj+vzBIEP69Sor8
IU8LIL+LdAr8CLjb7fynA8vlBwlpGAEnvBNZdaYa1c7yZ5EbZf3pJeRJwJQFum6F23RtA+DodMMT
Tw4TKvxLnsTRE4RlCwsayhHaDniQuMz184LsOhviM2OTYbi4WCQQX0e+FrDuVG3KkcOzRdioXc6p
t6U3wPVY01r9sS91pnB80c8rkQZ4lmj+iqxNNQwQO21Q9lTjCYBn1PZG1tG8zJlzpk9Kq3wJKFLH
8tsoQtrOl8hFOfYKEXG4Kc/npmA6wJ65bgGMrvmIU6h9SsxmkiHcV87P2ZDyKc8rwltICvVfN0AF
27HUXeuySY+Cb4lv5mpQ+hAEH1B3koB3GBxmrkArI7Lb28UFblHtMNZpjIpolZQiQi5yFeICU/Uo
o2Ek+ug/CaPGQDEAJk3Hjv0ZxHAPuOwG7VmMVppFzo5EpHlQEKq6K5WAtaSvE5kSHOMAyqGi3EHJ
Yb+pTOOKK0uSS7W1qCWi8uZoxE9BI9+tMA/VcR5KEh91ypAKCQ+MJ1pBsC/7jEySuRUJiNvSbvdD
Mc00uT6l7cmTzMHm+gZKtr3wNB14r9jG5Rz4i2+rwGov2cx2o1BKMEI7+dA0WzO9il0SrKKBtdlT
x76RZ+ohrLGpcmDVY0yqM2KPcrlXkHLzUtP61FMFMOCsLMYakwm/ahAG+pzORxAMq7hyhqiG040K
0f915r9KAKbD3WBDICe0EcthqOkR8LRSls8vi2gls/nXgy3XpVFIU7qs4dVD59B7ihoVNnvFlsBl
gNHPAajzVwYfGqMblChATjqzRcmXpMaACrCX7tFGgusDrDY8HmNFziC5F7HXVTBoKhRGxSTNboyj
5I1BXUCXitXqIsNYRN4QKOPnBTyL7VzSSzPZbPfdWP7oMXdj3iNvUT2Sva0BOQUhVfWKDfM+YTBA
vB3zgldtSYHkLdRpQw4fh9/4eJbvHMJpzcjkhl1Qjcmz0jgWTo9vxUhsftyegWqBmoAd+C+Zx1E8
h9zOAOpo8KloNMAEKkTdgg3RPQygVMJy6YG1EoCTmjmRshoMawV/JMXbTet4rkkBQO6WOXZIbPt4
dnz+3CqGPQtCuWLIeV9rAX9TeFeQYdh2zKvX2j0qGA276CFXmtcWVtQau7ZCAkNr39jCtMutvKtY
KcNua+x9iuUYIbrS5pPpTnUdVHur+dmIfdeqt6BL3wiXZzASsfZkfopcI/rRs0xtTj+kD8XLnnP8
I/+bdbRjKTbPuB5QfufBhNa5wVNWddEd4wgyDmv+KYV7kLFDjd3IB/UiCsjLUOen7NKeGzzYzpkQ
Mwj/4Z0ww/XAgxDGpxngtCO7Ra9V2Tr2cZhFiZd4+VQAN7mGs+rUaXwEqkh1RzE0+aO0BFdwXRTZ
jsxH+862hSqyrs79qI1zQshsgzc9ovDR+QuRcwhKvCug/mQn7Huh+dRBigHwpOliPxYQqAmXuj2P
SUIPGd/lOsitrAZiZHlfGTkymGFgBz1u+sPeNpw6fy4zhiC/rfzo4QSCB+8ujwrcOVSv5zisk+2x
t8IuLLo3F2lffClEyLJa9L1QR2zNcSMdfVSVzPl/S2o78aiXleB6YGPwHb/SRKTplbXt9Mk01C69
+jLZk3vJRL+mzt5SW/t1YYyqQgc58zgCk/O4Hq5/JrZgENk4x5wxmBp4ETzC15Q54WfpM7BAFIZn
luFe1UFmYE5CXy3M8bRI+Oyd76fIvn1XF0IWe5vmBOynQDj9czScOzoTARsU14kl4SpMVqGmFdc3
yvuxfJqTSUruEKlgf43I38kSYs/oVn/L4yvSBD8QUVNNYHOEAJ/qpnd15AuSZl3oYG7hiLLxfoqw
shKX65udI3LLc3uvnNDb/KgNkJeGNMHnEvL2imzTLGpkgMRr+utbvnJ4oVoq1sG7DaPHjIV/Bwzl
vZDlqfrpiMhiCYXiWc6QwSnlF4vv9MzB+KyhgWNMqApXuS6Jklzbou7ug83M7tu/g/nFtaeAeyfq
S4qFsZDygZBxNCWE0+rdZzxLa2JfepmncgFyId3nAkbttNDRUYiINYteoYtQkoKQf776tKnfqBYI
gQW1x/XltkisDnN0KOQovy2cHKrZtdk+Ycouu0TRVJyvu4ZMNBbl2K129LX1qk/s3KDNIgjRLn8+
gtEOwlOn00qC//1O2rpBGo8oGOWyUjioGVUDI1gNNuYUOHP0eV1hMkgh+aDAAyEOO1StNF5vb7Q1
fUovhStv2M1EdiwFNEuiLr+SRyYbAn/dO83W9VqQWqldtrtl8r88jwgUuGOMlX51OfL2PEhkfxvx
fpu6MDpYtSe4m/FAZr7jsxQEj9lbsW4e3DTTlKdxjzJ8uSJ/+ioMOOieRYejiY6BdyxEWTLHS3C2
+moxTyQKKwT0HZMNufq/N792KYmbawfQljYF1kLwla83uLM1VyXkzUnNrKeSsmSaUR6xXq2KwOoo
WSn+k+l9xBmS2ISShD9bLkHs9gOorqaJDKrvG3uVgTZ5LHxeAhpek+gOZV1LbvpCeup0lwg9kxoY
7lvs4KtOIo0YdHArpoOSdwHWU50CUkgIKwkzq5adHpRSDFzDTMzrcGwWfgNVlcpjAmc9ooPRBiZX
s8XnfH7DY9TAFFEfOz3EV2GHx5eTog9KE2kUPVC5QygmVdQ5GBkfDu6bQzaYpJzxHeODKo5MH5cX
NO3pz63wMEGzgyBSa3B6LgdK4JwTwfS2xbJ4qO6QTj4vy2jBBZpkLOr6AtvP9hcPxLDCMcpyma/4
okPspfF63ijwvSs3aU7oJzSLPOBRJ31vniRgkLoe4NU6ghCvJep4IE4VrmDSfk/zRcDfKkUUFxkj
ixnY0byAAHFu5BNXZc0ChjCaOG7HW9/sKYH6lq3cSPeJ8crCZOn89e3Eyxq1J1Jg6E5a5y1VQhyg
ASBgYvZvbDPnCVwcHXBqSuPkv7lx3rECmUXjiPcrrQAo7PCj4LR2/N263j1/iRDkJh8ArtMxuVgr
ms3t/voAtnEqjQsOC8dAdCvQU+q+DXmpmx3VVSha2ISBl7N9hrDjV1nipUWtPqKFZ0zMtfF6KLdA
8aIiQ6fgAV4Zw7JiNwXFfMDBEeiaGyjOyo+sAbyZSpDp26c1FR4rUkrWnJX+VZwFtfVjQit5G4wP
VPV5W3TMwaoWNT+jG5WbDCDY3BmuuzcGCDPxAaKbjtBqgZ2AKXnqcwXLii1pmENmf+m1aBcSEFn8
9yL3YXfxwmqs24Nw8WqLidib8cj4ioPdPxOAL/HJTLLdyPtLJe8lCml/3/v4zSIQFU6m12vIW57m
sbDSwd5zEB3gVLAASZEbtXi6AHYXY/nOrOcv5xeEYN8uDyZzxYBd0J49STut89ssA+SYLKlunAQN
+KtujlyVMUtsahWAfllGbNkQek9m1rJA9x/6VWtNNAUDVtfaCy+XhPJw2VKm2xIBBXlDnigw9Tqf
ohNr0aTtYPqg0/conmjVFHxZSXxugM4xoBFqSpHroMPHbHUwd9RZ5yeGRQvd21GHQ8FtDZTY65ED
WI6uSJpjiqqvulhy/QLZmXmJJqXUdn7n06VOGM5uSIf+ooqrhatrtxLvQ/o0W/mdHK04sXq2WFcP
GiqzWTDW7JXN/HX+Dv+d9NbXnNMCdmRs7DcO9iCIp1XhyopjmA2YftQLCdx2qZdXSWKkxHOhdjPI
SbnNaEPqv+rBLP+jAq/ulUDpP9zlscjCwiim29wlNL+TLh9jhyrDwrJmGBSzytqfGvk1dVaO+Pd9
bCwzIfH7H0M0YG20tnrRP1Imzlnai6WxT25vXRdK7fpSI2eUbx2jV5sTV3/q7T6JnIBxoMfH2usm
jjWWhdflvy18qAY+nNA3+u3ix756Gb9pNfYC62gdGNtaFzvb4dLP3jbqEMgIIkVJJz4RXgz1PPU/
V0llvTg0wxUl179Q3ZIVCC1jowENYEvHXIqD9TkmKDHB36uZJX+Yoj0Ct5ahs94Fu7dBKVVbmEt5
kFghx1z1FHX9NGuvZFHgTIGbIUKtEp/xORLbK6oQPTtmwPKLDbORqaT+SqaIvW6pF3Whl/zs5Wnl
XRbDIGqfOdL74UW13DXrO7qs3yKeMOPhs8UlnKpd5csaNN9SeShWxCJMzLqCAXQtG3krBb+b0LAQ
AvY8zEyAgOiX39itQXSSfPxbM62ugS9QNkR0513iTKbcRfTFdGJTJ7TZxHHFHAZ68fZhdNILLVEM
odHZnrt0szgBLmtaNTBZzjt/4GE0XK/bwVh9nm5YiKt8Jh+3xXUT4UUEHZ+jxcFL2KeBExtLpy+2
LtmynaoWDRHLTDaGPWupMGwyrHlO3KaVMppfgHEXxeXy8ZQFTWiuPTDQa7M/rXicO3/GqMQl/Tf4
FEd9RGMBVJwa6/UHMVwdxfGI9A4hbq+quSElaCqa42KfsjCyWw4C2da4ywwjfOmnHqr9mOCMcDja
JMF8FIKmFFcjmmtKtY3Pe7tzUOdJc7OQWC5iGvBoz+Z/+5Q6VNk/tEsuYa6H2cPQv3c60749edxj
RdLw0rE8FDKCXK7IgeGsu+Qw0SDTaELY15522ZEf/Y/kflZFq9r3q69Zu0LvNvtOZ4COdTLSkn90
E3HDdJvE4Vu2dDRlNrqXU9sXXFPOOT5T87BSyb1MTh1HUm7aNRjyXXQRBKuh7GOFMYrnL/dsmadJ
aFX8su9s4+sn5B6Q6C+htshnjCf05e6iascQK57i668Km/ff8r9hfvyRHVlt
`protect end_protected
