-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
03FoenT2QKaweyIjaeTOtUs43PyO0jY9YLGhoUuuQjFnDJYlBykZ+A8VkZ57N9SHOZ0mRLyhekRv
/TWxQuydnWe/NPMz6b4rC6nKpO4x4ep8UvfEpNl3ZQjMQhkxeTdfR1aD5b72XIK2QmMnZFOQnzqu
b4KHzv1YFKI07hPV0mCmCXwd/TKOPq5tngG3teJaBEfzeFm3Hg1vC52iEb5vf8wZJDr73hxDa95+
7RzWyXT7E3kR+DhlTsRN7Cypne1fangFWrxrEQYHsO1wz7XgVkMC+Ob1Oq0XCN8XubP6eLVHycPt
nB1uRljRi/2VYfiw76NRWEbPiz1k0FxWWbtcTA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13616)
`protect data_block
1UydQdu+PQt29YYGsfHkrUj8mwmFG9V95SLxRqdzYf77uBUD+Wq1uSj7KC2yEjNF8MfLEu0aikhN
GtGLbhIs7598Aa/hG+RuzlzK54cP78TegjPg0LZE6VFVSCt/DvpnUKBq2tx535uyIWXrbWYD4XKg
+nQSLM6TX2wDXXeFw/ywA6mBCFPk4Xkwx8latZlmZBWfeeAe8kubIU8Mldfu8M/34exkv7Y+yYyj
nawpaRTZCYSv90u0ByLmMx2pVz5+yDlQtNJUuGiQiDFNSvTpWXr0r3NeQSLrDHRJXfK6Y3UPOPrB
vdDUnszWOCGZhAGR56zUxGdGO6USCBTbdtfI9XzNBMDYG1A5D+TnL8PCXnwcKvsWw5bysjC6ObNR
1+Y7PLYE5X1SuJVdMJzW0fwvBECEowSLYPT9Uv3+Kt6SvUMBzyX8//msN63WUdxqfZFrzvOii/rF
QEjH3xI5F2yz84sTJ3ycYsdst1H7FPklpXjccPJQm6Z6MnvEr6fzlGIJ+G6SAQiwZOk+HFC0ROU1
QZ2dM9t9njR+JmUwy+auiN+H5stR86U7CvBVZps3EjRXPGC7l424WrvDEiv/CCEQnOdr3KScn1tb
2KzFbARWnUjNHRudPDeYhCNWdnSb+nZf//Lf3RJlIi9K7BbFELUtKV0HGHwRycsthUVRV6jKaZ7R
NGRCHpQU18QtcT/67JTpth9qGGTLB8edfiIDPNc/Lhbd+ttjUFc18+vIw3cTbOk7b2pLUtVgy41W
fZSZZ9+h1N1p0IY2v9C9FxIS30yERP/rki98HexamhzpN1SChSe66wTrYeQUqD1FV5OuK0M1YQjZ
D03q3jCC6CfKCEoa36cAFL7IkC+DvCbmExJCUbLkoli/9rUnNZ0UyxIxHHfZPtre2CrmYiR5TWUJ
JqDMYTp8Whwl5gcywxWvSIUrL970h0h+9yeZ5Mk8OTr/eM7YBw4qJuIF1ZCsrQjh6HlHE56hwUxF
edW+4/5QzmsGpGwXJMZR9U5D7nbzd1MLPgGQv+hj6NOzpIKCBZUSFAh2+g9kD2tt4i16qFhmG7gg
lffwqTSNUOb6tFVqeYh10/z2G7AVHUWE74jn+gfwxMTGXv8hansFW5JLThMgI7RFdLW+RZiPfd1U
w/VuusYe618eOU0O1ae/ZENSc7zXSWjRra3f3fDk4obfiNqO2YxA6s8CWIra4cNR4MFYKON0HXkv
cHnbiVl2jMnzLTCSSjdeKtZ3pMHIzZFM/odUKVzE2SBwb/bZRW2xIUqbAAOR27npmL3KbWylxVdU
qWQtj/+FFIdJdjjflUHV0YgPTvtfi9oa4G6uUK/++pwNnPtJtXBiDiZEN+ZEwd4CnemO8vs5Dy4t
PRVXMkznyBhMulei95Wqr77vrrI78VyIXMvhPrQYoTuuwg7Stipm4DwEAjDG81e01NYNtWhQu3DD
xl/xYmPW/gxvKwP1MV2VHR1SopY1tWKnrSeJnyc6LdA+CZywEC+lQckhy9QdaWqNMxV0Lci13Raz
gaYeERA3KzAlktfmQFoWyrFkDlwzAu5hR232ad8NBKWmH+lK3oyzQ3lkTJgU9/pd/hocRnUdSpO5
rbvELcbyGCdHWHYL4j41v5Zxx/L8DYPYl/bRzmYEkEFG9RbX0NCK5Aah3nTD7vpFlBPt+MGFFaNh
Cy2LLvLFVyNO2KyvgkZF3R/TzWFa+Q3/0Dw+VzpE1J9zinW5TF3ULeMtKQWC12yXpU7bj7rdMx5e
8et3M9T/V+Om8nBUBeJVwlXdHwsHNVpi69TTalCsGg7eD5f7P0KL/von4ymGVqXp9THu2cflwuuL
Is93rBbSJyFS8SZ+Y2QfCj9sGkfHdUiAPbxB6FkB3JDZAttPU6mG+rPq4+B2xdJuXcU54GzF/2qN
L6z51qcNDDr1GShBMezJcAoRFb0bitPVrl6mKU4Bl6vg8LBugldAyDrg59D5hU4G+Qr0UKwWppQE
eGjHquucuouHjrUdGWR67mO2C/BFblqEUu/NFinj0u3Kg9oE5g3mj+8KTCx5Z7SaUNAfzinE1J3I
1Qt4T5DO269JcE0XPYG5BN10w7qmK4k8nEztUHsbBpJmzTxJ98vlJ2CZtGhcgSAigPP7qYXaSSx9
RZVFicfeoHPzw3NMydyrHNXr4m+kSutmk24xRBmBQZ25dKRFMkZHeZe561k7jU+OS34noPGWS/g9
kw9vwYDE4HdRtB/xsEUcRfzef7JIwB64IdcK7Zi0SFQVmVusTsRuGqGZwzNQlmgDbGf7UPWp3nj7
J1Lb2KREU1ZrK2JxCazG8kwZ7y/0gipy+4u8XbikbOmkNeNAPJmgAHtUiZHnHrj7aD0wMJZZbovC
wke3NjKYxym2iXdpWEQWIll1+IjMm0ZTcKGFiJS/DD43utoRjRbyOyFZHHwY6riE80GjustjfTqe
hMuOZjyl2J70pJIaKkcJLoNtgGjqOHTIX2n7sWnE/dvEZA28RVgHqI3zWczK9kN0SR3vCJlARisW
Qp0bcLTKDEUDL+H7D1ht/gCReJk66p1vDVAX2qrmRXyC7zHUWCspoNVEFycymKnXwTr2hXlkzg0d
A+5NKDgibD0cm3eLmApFG09pEdrTEMkTt8d4ODDrC9V8JPbh8nor3oTEplkvAPSJ/yMGmBL67hFd
WPoWeV1RXYOsJlbSfAOwHHJJuiQd4TFxtcFYa3VFwF0Z73o32ffLTC6e2mEwgXuIgwEchfSqQ6BF
lExU84ejV3mz83k+cz3qyH4vHYlkdpLB6groJG0oIVgGvFIM/36FHSlc8SNqeUVCGMqGS57kvsek
5uRA16GNklZcXJzhZ5AFHWXAGdBhGKLJ8JjFDKck4QjY3p9Eo+KFSdznFvugHXV3TzHZ7fADpe5E
h/cMrMv19YNDBuHQHIjsafbMknI0cvGLStMIybQ2FepY2/5DinpdEJqYnr3hD/tRIyr96VTxYvYr
xariS1uOGchfad5vKGwZ3t4UDv6CnWOhteGUhJ2F+lc5KqBl3KiuzmxhI9xUtYpphXHyfaRw6PLT
ZwkB9oMh3XGRf5jdmnZupj2YpdKmq0VwY72NYMBiY8PWDRKovzfBqMn1By7RMgZCMFvvUJFhnHwL
pREsX8+NSCAkoqEae1CMtPWjJeQS2AXuauN72SJEFvmUdRpyg+Slnbv4Sha5bYpMmOM5PynsDdSX
aXDnhv2Bq1Lz8lnuvbYGAjZ1zqbPvKqy3kePm+hfucLq5dMcGTYGsvuGCsK/O0yddBAcwpQ+lv4G
TP7Wpg2q1N5TbbUMZ/0ljqBhwuHy7BGousIg6vGPNJ9N7x6+56uu5l8jFvw0oK7KkpDUIgHK9Zcq
lUUMl3rlxSuVbYicipJGGx/mxnd0LXPjAAlZFujWdvT8tM+S1PUAlb0el1pcLxKeKh+eK825yauR
Tie3WfJ0ClLzFasDDJWMNeM9zYLyxIqd1VzQv+Drtg2eVSXwanD8uv4pKe+iIYEMMVEq2YlKdrje
FR6WuXCagsmenU9nnJkKw7zEGV+d4Ucpa/GW80O7AxVVHGr7XKN+tn5XW8Frjkt8OwwKb41MLbho
8Bj7vJakLpjZwFFjQIh5VWIvLv0rxqXUxeQnPQ0p7wD0j/vnAy9LAt9Hij+WA1HK2bZqHa1NKlNx
3+a3Eksb5fQd1UvAyq4MKmZ7SHUQ2oPUXhKdQO9jX6wt99xVH4QKYyggzszPr6jzUykxVmiSuWUd
v4/zxaHjcZD/HGtg9DYyy6dHa1mpFpyAMW079oGZJesFDiX7Z5G9X4dDpyGY6GpBXIpfiDE3ivPb
BKle8pNfX6Tc0fRfibHdGYxdiErWYze8bcx/4033OFwoQiRufoHiaWeCd3GAsqKZZusxW2+xL7qd
WohGfiqKCohJGffJwYySrNMqxMwLDwpBe/Vtgjt/JNP15d7Alb7O8zi+thEo82oL11qTpZJGUemF
ai8vvaC3QtsZpql6/Lg1WfkDc++MUQsYFnW11/ka9exK415OB6RBxxKIzzz+x27+Y+yl23lH0104
jV6S8hOrt+i9lCOOpDGVk7SI+ldrJSYFi2XESnRKTZXRxo0P9nVV4lKbVcBj7uz31TsxGunRmuCX
cS/bfyYPRhulc/EL4pRNdVi1EJ2fPW9W4K05EbCH1gluVJGE/ErMJcwMVFn5xSSJlUJwkJW7xQ19
urhJ1kItxXW19CVktW6kII11HqKpvMTTCCBaSmqXFFtwgFXmNhqwXluwQxe/Y8iH3FslyBg0Lql0
7Baej4C1QzwlzDHi1+JxUwrS85+3mThZvXClebyoZbfXjptof+eBP4DsferkOX4wtOF2rBGENEpT
Sd8/woqq/GWT2f8+2ZM4iWD8UZyzeyInebZ55gJrqZAb/4myGSnagzg5u313GXibjDveTF8LB28S
eLdZg66GG5KLVrUHhJUjJiDvS2WFP7NcouI5ZhO2GRgLghAL2g+p7428WbMLtFDRh9yE243UQ+eE
3CNBOsYNMJhzHr94wle3sGLAHG261X8asUW09rHsmUL1s5McGU4csHRLd9CBYvgNcMItvorxHoph
tudf5/HXmY+ICMKdFC86BGzfydpClfvTPqOCAucw5YkPA5WIn4o52k/nsrHkX2co9TD+4Bw8hDls
7uv/wwiFMXI/qRoi0AE0RY9cZnG/t50RgF1bwc6Fa4J8Hh24+0jlcgTXc0Gyqfo/YBOpRz5wkvcs
fPPsBJbeRoBirtIaGptuFE65AHLkqRaUAk/eLloH/PPFpQ+ktfV+VL12+b7AK4VGDGDPaKyUJOyQ
rzei/ECvgZax5j6qU5eDJldDmM86FpAsGsAzh2dd+PYZwhm8M+8kUyXA96WjhJnob2P6WS+4uUvn
poQlebMjDfLzWdWNGXmrrdhvzxZvfO91frTqnTX/rctLIkYV6vxmRKdRl2a9D4WWz9gFDD9yqc3/
GFnsLAafwTnKAgOzpVmk+fd8p4d2mdwmhk5im2Akd1LihplT5a80PeHDxSb2sxvW6ME0RmSjM27k
YxOSsgnX8yHd6Rw+MO+//y183eT2ZReC1/zMqJ1fvLGtu/YGaomuwlWsvkmtf6YVSVOw8bTt058e
qq9gNsNZGxLgELuN/YutyQ6XPOF1h/yEiH3fQx2+762oQqdh8vzAu+xe2uhx0MXL0aJEKxa83iMk
nv5LEuoFDuB0O23vnyXyCwvTcjy5BSf/hX/JZSWbEvb3fQJiD2vZF+JUzx3iIaexlDRC26fc+IIH
G60wd5h7J/AF3+ZJzLt7YZAVjtL1yJFw1gP/gsBQXYUDcA6Un4qvNkqzRYElfvs1R6HzVhCwFPCA
NsqzYCLMuUpu4ze+SFuDamBcHAfVwxkvBpWcOHIgBqGrEsDNILiVKFDvQmcclx4CxeY7u4UHdlLb
SfwZH7nRqq6XsoxWSJvUUyU0ymP90lKkl1j9Pes6ZvQb6NxOE0hWxB4mF821tDn1D84rEJGUeb2M
DDm7GCRDfx5InG17MqnCLW7vaqbTOzg9+IkJ/w4yscPCbC0LI1HwmVh4NlJ9pbywoAlmb9h7spqy
cstEbzlUd7HIYV3O+uQg43CjxTqUZryDR0wiYTIuQpG41jbOsCLKj77PiyIYXv40RAW8epCq9GD8
/GX6981Po3xnsnxLmJrBWXLDRpomGc940iL2meSze3f/YDBB9ssnQ4Fpg9B6tiJsrzab4PvpNrVT
uthG5Vhxyfl0FANWQ08xZW98xeYAktVtZPymgwVbvcV4GoN/RUMmjHpBzh169AIKgeTrirBKTnCv
nNkbgbbV35zLNyrdLtCqtWg59tPH+348vtcxkARLr+UhpUPVg5BuRPmlihjXoJjm6NTGaZr3XmKo
GWPn5gQhkE5dJHkzaeqLY7xjCvWrv3HQns61E1U/ja/gedh4+jdUAwLedHNrrgmx7jp5U9BTUmHW
48+ildFX0Sd2utQDAbnuO5djJIY6TX4aWD5dODG4ay6AMOVy0L2ZcAH4Kyf8lrRvo/gKZNsK/aIq
wLS9kaGHNaF5XZXBhsZ2xyPkXyUewtpzQPBBAvB9zdg1fBnLFtQWzLEbVIxwiMJzAhSyp2Neyzqh
TPvOwBYj/j4omIs5Dn8PuW4i5WioGcSotZ8PkLiO3mHO/e/8WkUFG1UTAgarJ3gn16c0jWUYDJ2k
JAD0ffvdY4UcIG0MYKNHrWvUXbOPxN+lB17ARUspu9w/dQC8HYrXuUetBRFvmSLJDoW9oNnhUo/0
uoGeK4l5O2nU8sN49tYRSJq6gThYjY7p1T1FeWJ7u6bu7TwTwEr0YsYTmjDnRyOYKkP6G0v8AYeV
FB1bulESs31WR0426qz3JLNDzjHhertpsxKsmZlNZU90v8T0UbduYEmvzzzsVNkSnNSlAVpF+sD3
jO4ueWNpoyGf3Dhh2Xt/2VVCyiBI5vqIvlE2zBY77X8QMHlse/Cl6CeE/O6a3sRmTIdKW85PU0ha
Sc94VUSPnfKtqEApfFoQsPZJ7dEDNdNIar7/fuofV9bwGkC/9ut788hsN1ViVprgiozrMNGKT0zB
9sJs/qwjmcs35iBAsduNfBsLxtCqss4hkxiTqWpoBKVPuI38PPqHjbqyUzwJ8iDFDj/RsDFW7WWy
aVzNUKImVVn/hglrmkZMTLhTfynPorrtbu0WwbdCXqD2+UZ/qC3TAG5F+gLw+YGkijQKj8ecBic+
WJRKHqZJJbTxnhhI7hoWPmDCD0I5h0h+FLEnA8PvaiHsKurRy9oMLjI3thoBOqBkgdOvjQIwj+A7
hM3g9D8YpTOalGC55oA5wjfnqK9w76DcK70Kzfbs+o/8XjZkq9z8boVqPiJ33QTU45jqVJCnBvqo
YdCt6c54tycGsxNEVbqr7sVmNZjrAFYtHMqNGzNDRD7I/Go4yjE6Rdb+gnrHCtEjUwHdyCVnUaVf
njVzKscTij7A9H+57YFfWUdXik5KNlHd53PH4oCK9RruF/u/iDT0LgNXQWqebV2deFpqAWF3d40k
AMTUBKcnzhC5L0fhSSJdDNjOYY0Pycd2N9alkmULgA4eywa+2zsx0wYSVZLAtq0Hg2dUZXFizL6y
CjzEBHGBitx29fNOpB26rQuSr91Y2boridrqEU5ZXzlmh+iTdtMXIiOSbZBaFVYjkiqaiJHAmnGH
MJbpq4+vpQF7kMbNMT54o9GOej3LD5kluXPVS2okyQbX9BbVV7DrvD6to9VdRCAnBMml/CjSZmey
3vl20yESxmaZs2UgL7iXWpccGKCm4vNw5BE2BGdcdfWqAC/uwfmEvyyTkf5mq7O0pnQSSk1HczCK
X5d/imRAR5oeAIkmkbWGZC2c2Zfzt6o6jZEbZ/sB/mmALW4oet69cBYXMYjXbJVF8Ru+t6MvTNVg
nwlUHH0M5IxGZrVV5oYWAQrIUzGqA17UGnW9jwuVngpIanvHtNh0Gq6mPV7qGoPYzzLcIjyZrKix
fJ0T6BiI41Dvbl5/9jbzfG/b01oxObzPyovaVpMpiZftnbnr+65IferEY0YsExkvUy4H/+T3UpnW
AP6wg9NQ0MOb/AFrAkuRpz7FkIZRTzB4Z6xIgXcKwwaQYMoPLyw9vBZCTokTcpn1pAhqGQZJGX0e
tJ8ZBf4d0A7fpAZksOLU3GDN3Ab3quNsnUqLt8uH35VmokaNaNTOxePcTOgMg6haymnHljjnb0YH
9W1pbRSmG8aMN6qu/PtxnDyXzr0xhfOCjKO5c2WsIGF1GWl9AtFmpfeJNkkOTVaItVU5GxRvlFZ8
YywLoaIe+USE1zeEq3oTvAsKUnpf8Wot+iBsbmXHcS9Iarwv4QU47e7DTvUQygIFd8NEVgrmBLzq
uPe+wvudCKu92ckXivBVD6sN31kgO6hblbShT3Vo9dRxMvvEFZzvzxffxnyHuZKIYp3WfkRdVBS3
DuYeOIfQN7n3Q029PYijJWPe+R4Mg5ub/fE485G70Ugfq387KwY5F4O4ObYu5X1nAzacdHd7dX2I
KUWhDarK2JLTig7N1daEF4HaCPLXvzFoFyr8U0xu7ROYbx0P1SRjSelM8L6dqH8mLLXD7rrKAaRX
buQLrwzpSWymFWlsaLholP4kEBGhwkM3Dw/ybeZwL5fYwyMjpwmTgxtVMd1JOZAJM1buxrlij4Nc
KCj5mxGtpPuFrXx60RKhSg5PPeYt9kckcxf0QtVj0bwAEDAni8k23Gtr11t2bCjSmO6LDcC25zpa
dLuVqF46594oXRzm8L4H9sPOm4E6fgiEhywxMj5aR1ZcCHbwqbTTfQ5IprGmrpcAUQatVpnb3Lig
hUo5MYXlrxQfOnk9irvJg/T4NriFL4ZFzj25+b61zQDD3F4FBUgfoXZPVYE4Aobvl0XvPq1PSXOQ
PaHxx37Y9TAGI0Me/OG5Ek8TTIXx+9COUMaX6I+zVLTN8gc4+5ne+9xgvQdVseIoFtlaN/F3n3Zj
SSVzheRwJjOaO+e8RqMKpJv+sSuAhdKqTi0yk52au4T7AFZKwY3Nc3bIBABDij0cNkkCrQm5aILF
MvJjq5Jvt5SLP1r/5oaMvTGJv+h/xoFveHdYh3fNueORKnxxhQkwPS3gquy+Qlq3onUaVAaG/omA
eK9dPRZuy7H+gW4MqFEocBfyaGYt/C7N6azwV3LDOWsMMhxynOwlZyd8stn/OjQtkA/1GZH+HQIO
2HgoHZBXGmCzWSDAIJewaLeHzRdFM6+hov6YYIdLHfbZ8esGg4DPch77cC/gkk4imEzxZuderzBO
8sUIdVnO40BoHlw3wtsCBdosd69NK7NVuuOvjSfPWOcGqqFDUq+If2CC2DJXpJs0ENEo5D2eCwhU
gXT4wral+p2HsSo9ESztI1eA+mdQeL6NOV1gRMpIa2p2a2mL6sPo1LlKS+FCsfjyrkG7Puawvxyi
7oG3Jfb/bTOlwPc89x//azxI87X/3PusgWvxFEVP/Ruq21nS+7JkN+ji5IciKxiE0XsPyJIDkKQS
hajWxb/BJpMP5ul90jBHjJqLSB1EsFkqJ7zKtGRI0B3STfQJYn6XSLtAqYw5qXoLKWxr6jUXF0mr
ReKS5o/+PxbVeJENueChKsek0zq+QxXIGGwClMIcllv098OeG4EAauerSHUIIN/+wld1i3eqsNZY
ahw47ejdVuD89OvcQbxTM646rhlnucU7Gt3Xu6zQz6jPtIUBFD931rIpT7SuQNQ/6IMgxhaECp/B
EWpckt05MGECVSZnvSn2dIjEUywNRvIOeTu3KkYBkP/RO86z/sO22Y/WJxB5tENLh+vwMENrse37
ZKJGAXQIFPXWaw8snhH3DrA8Z4Y3arPpmkw5xGStRw4KIGH+vn+jMySWwYB87QR3kASzGiRSWcx7
p04VuH/WmBhwAzgv1OoamdFza/vNiTvDlDcvS6SOfjqFnRGu6WOOGhd/zMZfxXApMWt1TreONsS3
UrDHkE0bmCRB2MQ1rf+Eom9gSFn5Q9wEIhT95wC/mAxFplmXCRoN/u5fWohHozxRSE9u2bnk0WFH
zqU7e8ZLNacuHBY8sKSDFJFqU/WDfZ8QprPAgwBM/NCHkZXrziUcfKbQh+8AvhgKrbmpHSM4+bho
WsTQwLrC2v6TjjZC+E0vIcRuNw9ccQs6xa0iRwFx5FUIqo+K/dnu8DgfBGealIiVdMkX4rcBKov0
7OLGXAEPYA/mD+JJg8pfAx+xA5HlfVTjWch3QIjlnKmABZzjFvfJl2EAY4D4KHvRoB+CVwHfrPrA
7Rp4aeYGuWLmxlP4lFCi5v+GtiEHIBoGPygoJK1iKhlzqR89gpPIb5TkzOjmCZhRArwcdj69KRG1
UmhnJGneVQMg7hxomLHdSENQR5ECk6ZMcOYpGzoOo2AnMMZ9pPMiHgZN/eInkJZxO20KtCY3mYAb
2tjA/4cH44Z9kx6Fs0/QF4wc2jKTA1/hStLcPBI/MWokOPD4k5n8Y52Y0N5FFtk+aZcsIdjsv1B2
+0lCId6qU7qMrEjt5Cn4tCyLF9AhECThBHkUmdEkbpNktykizIMQIf24bJMjgrvs8d1DzP1FKMmi
tt+jrlXlOzOHl0RhVWaKu9ZMfgFZxExR63G9fartCd7BM4J8jTLCtm60Q6yQjSSRX/c35jYQXVxc
Hvw/kawLyjoL04J+9mh0JUCFWk4cCqVHqmPQmR0ohWszX3T/RhSCQ80aZIGidtOxn+71Rz9LVROn
tgu/dC9iheVjobXrFJpLoh7gSftSe+Wp1CT8sRUbGIXrbppa2yblYlP+T12kwiwsQY/5RpGYtDyc
BVSLSAvsOmCWevDhB6ZD35+5okSEmDQ2C3hIragudbnwuUEdzBIhACBo6mDgW64HWEM1UZtqdFsu
KtrCroUzYnvyQK1RsyjN5UPhBzIevzmvN76zG7X5xBsFWStQUWJMj7u7rttlyeICbCYNrJ+AjpTM
xrFgsihshvXGzxaney4Ik+gEgEMGVyrb2gfbcAzpzhS8uPZVRjJ53Qs6QSvGGhmj89LG1U8wPqKK
iVLegUAAhrVyvqprHZyAwtQkDB8H4PsO7oKrPsqRBN4usvkAGF12uyw2WHZ90uB8rc+nFZKgeL5C
OXHh2mz/tf2oSCVYFfUduULueREit5Dh7L9bOM/BN4DxcNQcS4RCbkhbJdp/9lqKuBYcgDOZ1yis
3Ku3aoGVh66C45zWfz23SRpPwTMcBZGzSVvPqF3+++31ToEjDHV55MKsp2xMfc4Tj3V3AU1829C5
dNdNh7JYvpnsKvqtDchxQG81W0egLAocFcxIJRer6Ox7TUdlmIa+qfjXp51qgXEGDRV6lRq7rvtw
gDUDYWnb6F4TPJA5uZvOO1Dc9E5DbGMZCRTsN9WlQ2d5VJR7OfxeykDu/XeLAtWtWgGakNUDHRSt
/qoS3kcpDJTDP/pjCg1dXazXlWt6JvHfE48AR4g5B8DjFGpeZg2WMhnWvP6apIG+u6wjodDeZpSV
EReI2RC6H7ArxlZcdaEeGEc85GY7Ufe1hLcflgCfITeScpBxpUWvjZiSYVd4T5kL6mnrrNPyeccz
5pighhz2Jibql/nawk9QLTIS7Uy+NZAS/iY4BlYBFuQaM3mt0Q89WlT8McdlyeXhOrU6U+UL6K2O
Q8EY52iQtknAAESTO+IEBv7k3KVra1sbnTSBO6Pj3FAQnEPrmkW2GdDGlsudxlOcM3wtH6CbcPXO
ACRONfBSCe9hXuI0QnrVKAyubvVK/OqnAuHIbp3ZqLj4c+Q71v0z53AsblZliDlPqLiF2OwS9GZm
8W2fZyfgPPxm6mbDPOtFaw8u2Hpljq3mqJ1o4j0HRYaNdGGC04qL9qvNeM8j5dLkRiMo6u+W0akX
qKac60HWTIUkdZu/1DeN2j8L/R/jHiq0SzP67GeFrzfR9VYhWlDwtZrPw3mhCfYHKmRho/t+PeZK
TE0bdYlkXA/HS7JsgdqsYClALx1Al8l9zlvX3JKcARZlM+RAxuUJ9LNCQZbvluGKQLPNG+UzxYUq
VS+FNmo5GSUru6ho9Us3ygSptNtrocJgioPR9AINI/7sP7DBwlsfmm0RTvdptAUshd55HG30SoMA
IFU/c3sg92L8YQrHsCq/zm/c24Zc3KPSE4n8NSjhovMeVNd358iKEn7B+e7wATTUXm2koxv0GJMe
tT95q8wEn05dAlfxujlQqpl0nkcZyr4Vqycr88Lic2hf66zs2tSKwTTupc/H/MFRMRmdiseR8EYM
X7v8w3S5tS8GzNqbT1fhhoq5hR4PvWGbGn+o2M0Yk7CkwwOQ2w7nokKiWunuYcEl3B7g52MmU1tZ
LUUZj+y/Aue0QRuMbdFjHYUTsJ5gh2yc6e/sl5uaGGufclnnVG8dyiExQl4MXaKlpGkIW++g0Mip
8dNJRNBSLqgt6mAXTCP6b5OYBGKJIzoENKLYq/SMhUcQC9BQIdm01xcYstlrXYz11ihxKn2XgRBb
3cNmkr3w0oR4b9CSivpdaiAnm01rRzt/T8FoTQ3Nz+ezfEAed+e59IaXQ3CNz5aTFHCxwLOGaYuy
w7nuhGC+A1AYu+U3q2rX1ma/1ICdwF8XdQ1mg+XBGzjE0/6VChLgYJflaWFOhzZLJ76UGXZ8tVQ5
LCldRudS6CYnFAAV6vBznhMlfCBC5vTs1y/luSLpzEdHYV28ijtfGmL6gkjeNgGOTdvxjvK33VPW
1vtkGTvQVmf3vqMxM+H8t2+CbZY7V2GG6e8xB1AMK1XC5hGYuck/ymKrUArONgo2UDdzcFuPFm45
u+vSLqfsRCdeLPUWmh0uiKUy7ik4SlOmL+K4NIkLt5CRlug8Ywnd1HO7pdsFIOaoPyXu3Uo6sMAx
0aP2caXsE7bCiG9Xw5v2MoMJ+q//Lmd6IhqPof9D6X0lv5yTNIlAEC5ZU0TCQfcX9mgH5QMPXP4U
JFDOliwowvVCf93mq4BsWuCpw/z0E/GUA823KoGgiXtyT4aLZaT38UihD2Z7jtnvksXEXtAkDlA3
fRvv2/SWdJWmsmz7d54LCxqzeiqJNKdlA2lpoglXMPgeMTtItd8zjiAxxBb8s8JZMXDuAIBATZKy
ZEg4kpr1vfHP96G/GTDYDZjeY1wsENwRi9rdn7ptFiyaHGVMW2A8OnZ+yB6da3Fy6FvHH+lwZTUi
t2b6GcXD5Jnyq9edi+B+ZjgpRWHdwYlMfyqqS3WuircROxNhCAijkLr2aMix6ANW6vEmP9LKacKs
GA5PNwgPxCYyGqY7rSJAmf+F47/rU84+0zPi4++pm60E+g7PvyCjAoikxk5Hl2IQA0wK1gnKQGI9
roVsSJniEohHmwyzeM/nMKBzPsJR1P6KRHlpOxSnDTB0Sy5ovKRYZIeOfzGBQgLEs6Qr1tSgCVyR
18BswOcD2IkXYUOsDJ3AH/FvT3BNeVJcHZwENnBmsfesF0vRAWObjPWI5TuLgvl0Vm/zVN6rjYEF
snBY7jPGfJVt1M3/kpwSytzAt8OydBR5tBWqeow3mTxLT2A0mCcvvtTAJZo6Tzx9d+xZa0fGxTnJ
o4EjByFHHtull1Uhfi/EpzJVh5rPMko0FZBrO9xIgTAux039pkGEwC255P0ulnpqsMpKiTkDvDnx
cSephDEuJHkLCyePEUzmLiAZHAN6FtH6OpS2WqJ+Xy5l4Xou/cV/n2b6VCAlKMQpTdwS57v+EhxF
Me3E7vXaftF0ZvDFa0oVKddh7i/AFhBw7t2XEceNst3DOIpq3w51Q8zAU1wOcfRS7OopYbmb+BVA
Ea1dBoVk2oprlw8PN1NYPMg0xKG5QfMMBKffQUa4PuBgHfMvwglK6ty9M8RK83/IDEtShXKwwM6S
EURKeilO0ItMcryciSRssuyaX2oGQ5Hb83P/p6LqkmPOP5/ZG4wtwdh/MJ3Qr5yroksZ3DiNV6+n
TYLZ2HoEdebBKO5hVAnUdmdtqL6R6xs6WtCF6mvraKDy4YJTQchXhnbLwKu5kI1NpVasOFzEg6XS
GEILMOGGY53/2eLctzgS21nBW7EDlmd/AamY2/KtHevVrsc953zTjMWeeahAC6rQWGTAACTetYwl
Xi8BMQzjuNhz8S/aqUj36JbRQL9j3W+QX7mrSDhWCJODUN9qI3x9EbHjNGzM7bEN3Za5FjBEshl+
7EaYytLTSJw84Dfrl7OifGtbEyOzkCqOCgh6MS2H8uKRSRLadGPy1yc63Y+eR7Tp6zEhVZR4NOAK
IaQKRmQc1Ih1Dn5Scd8p8QDWAewV5lVUM+LGTkhxhBvksalL51KFiUYQwhbMUOoclLB6erpcvd5H
aRR8xGQPS4aQa9mI6WHXuukXJOxDGF0wz+Ct9bzWSNSyvyyNtHTC0joJDS+Mk4/QQHlFOpy4M01U
xoEJ1WxS0YcWJKL4/8F7vJXWFDq8cN1lMOJsxSN1wBKmTvMuoe+LcLYK+A3j8Y0spxJ3xjA4OuXq
Bn5IvECvR/H6qNeMB1ZbuOe9RJCXg4Ech2tUxvkaKkqJRik8RJF6qc1EZYUucKQeRdVaU4t0uRgk
o4xq9qzTMIfYoHbePXoQcinxj4CkT8dTZmkwGFlH1XuWc0Kd01jYToaSoizclChTOUE4qhqOLCKA
IwgksJw2pfUxnxajveD0DXUuG0WJungwtbKkElDh7wTX+3kgUXR4SyimUD9qhcjshQQYN9slm6Rd
NgBGb3Dy8aIlmsRzzVyQLLVPA0fQ84xMCY4Qj2UR392jySVf3umLDmQQE8QSroj0ndpUWBCmUJxH
eZT85tmMtY42f7Z69DFym2kQPMvyakzSslFQxnRy4wEvEUH6LV9xad4uUBjtIpAqySXTCCOYE7dK
b4ilV7nU/kTpMTa4pnjVSy5Ttma3CUk9rzLfXxMpk18SgCf3ofE4bnlWKPsgrxNDxoSRv0seiOGa
/MfW6ZLTGV5I96aCnuDH8hEtOzay9Ak2B4MsnN9KW0iWrpbNtsH5Pnr9sU5YJxel0CUBpJS2fK8U
JSxjDaUjKlzzhUkzENaCDqv5wACCJN32fXSlpMMW6PH5uH/egfVlqiUnb9Uz8vA7vQj0LM4rlQTA
lQfhFP404oAahB+uDdBWAd7Hka6KMRLbepYFaIJYVKdlcAHaUHBIH8Gkmor7gB3KoIWsNt8mB3I9
UiELBtf6kGwjl0alM3WQr12/48MihuyOMWT1SyKDQs94IabCVtwCTX6Zo4D+Rb6virzuPD9xl044
8FdLVSPdBXG7HP0p8GxuVFFK59gMGYqMRL+BHPu8pLb9faWeLb+Xt4VryWxITca44LcJKBXiAQGm
QuoKuET6CScmO6dS0PlxwFb2kja8jc9Vj3QMZ0VheWjKxlLvAe/Rc/Op92M+uTJQE9AqolAFq3/Q
/sAXy74qjXs9hfWwqkqYwpzDWG0B2neVqnMDcgWE6OJp6Su1UA48Undk0OKRVHg/emaYpqPqoth+
G+h7XmJPCssu++fcgWDpZ/zY5hsZuymvtH8A6Oedo+VspBo2pDpahxC36PkibheOng2WoakMYNRq
MMV44fUxROq4+Rge1MyiITPqPD24Pa64R8HD22CoHUjZxGhu1KaVLuI9Y2jdq4L0aP13qCYl6oUt
BExM83ZMvA147MLe/LY4Hh0JX+Jdsb8ZaATYSAnlklN276Ov2hGG62K4eDw6d85MIzrntjOqS7Qc
nTpfmPkRFgbgaJb08m/J+PL1MhUwt5AmBy2NkijU2HuMVap59A1zr9+scCPAVPIEG7uIfkxAWX/w
irrLMLJ6pxPjoUNo/b+dEderzkGSV0wD5UzhSlGNOjfOVfBEcQSzrsapav/o9rywMl/8Fs+y+g9h
Eibi5ATGQo7afHz7zyyicEZrgGqQfOUiaJuee8YSQs3iMYde+HA/tpHyQnfxEToPksnqT0jtjS/u
jyLp9+gv5rQertLuK6Ql/CQ65vz2vw1Y1avGmmf7/9oDBBu8ZpSmHAAz+qaPBwtFCIeylgIb0lFe
mZfAdXzJmUiU+axvF2nlM0p1gjaP2CV9pSg91PF76B3sOl41VmGaBMW0APC4kgCdaQylNNMVf/3j
/ictu8ifEzsjnts2gJ/d91pZ+CzYHEQUTddKbjJlKXrAvwmMs+WSbT5/v1o8710msH7gLBs+2n0e
ADz99mzfuZ2XWoZ6IHhj7G848LwAOAt9Zx82yCObR6p0kHK536X5F7D7FH4/pYjLyW25a60RGekj
7oGV82NipOeSRQVvftne5azmxEcgFV8pRWckKpEClSU6baPwO/4OwO8mpA2Ygi4FF5scxOIQ0ESs
4SQXOQ8zWhtgwe7g6YJdiNO/YW0OBaKtbWGHRXYdoyDMX9CKe0rX6fbQZotaY76qxnnxVtmJtd8n
7tKW7pgdpleqLcBKZPthz5rjqOvCi4UleJqCkpWGIBBPpjk/hyZw24mTJsRG84XSTSYPv2Epljzl
cmSjJTNgBCVHqmQnThMbW+ReN4vRWvkPGq4T0K7v6v08wGSwYS4YFY3lGsr3xPm1ooppH+sopUUZ
mmYnXJmGSwmN/j7meXpaD4b3SISN1aRluiaBvQH30UdSR9jvHj3QFysCBaIT/c0MQTd4V4JwlWAm
Zea5/gSvkR/Gvt2qjlJaxltd8hhVDX32ZA7zjQqyLtEc4je0ipU+IJvPl9fUBPEwmdWnVDkExAV7
izNcZhg2ZasyPfAen1crxrr0yepyEDR2VoBJSojFpuCXESiQm5szcPBHEAXVKULgfssDAQ4W466C
8jCUcZ15hd+KpZbcu9IEnWtOc0c85Icz9grIbqu5nPZXI7IqfgFtJzsIdKBkV0Fd366bNMzLjHEK
Pv4tU3i57ukuSKLAzRR6N2W/jhfQfTT1eeGac9wKa4ul+UWePpNuVupN7oBo2J+HxOwQoS7VHc1e
RfeVzwkpi8fVuAHFPJFYyXc12JBUfME5JGcbNAvusGDGOWbmxedikwSe4w4vtWzxFbvG/Rvweeew
k2p3z+hVcXfMtSXs9t4gI6KiTkbyjkftjhlq11+/hCuwRWjSiDumF5ROX9vPZ5D8TZxukNzzLcLH
3f5N2SoDX4Q1h4eW+63ntd336faW01Lks1YBEhW2Svjy2B0DGrlvIyKxV/nRAW8w78ncFqH7/mM0
NB0jK+ON8UDxCfIgLU+Cg0X6GkBVndTX1I+zQa0cCdVyPap23r8XQFAurWZR7+TNcVxCVWuufk00
CqbFnyfGGMjPA0cw+2pPC7x/bdX1LU/wHXv1sFWkm1DILOk5ZEMgMcsfV4E4luODh0ykwmtVbRqu
36qlXv2txjUqJTeFUGwR0OAOF3hBHBKQN79svEVJM9RFp6FvkX+2U2gx4kf6UsbtS1TE9axIOOgK
DqCxj7z7KQ7tqQr1IS49AcFjiQQu0xS3ET+hYNDCOQrpsVtFSSI3CZHaA19Cf8CFSCyS5nD/uDNz
LaTHxAm2mcCOtV/+GPnoeGsf0HzafDbYyvz4H1SMJFuZVq2E5saL85VYn+D+a2T8kRsco474ljF0
2Gj+w3Fb19Ihl00WCQiBUBv6a5Qmg2UgrIPrWEypNsBd25YGYVg52+rfOfujhoJKuzTeGU3uVyab
wCpJSjSxmiPN2+sc846JV27c5eSMLGqpnbxOH/MzGBpSoPGlMHEAmU75xkEdExUsnlsBMtx0B70q
LOmAVX3N9SpLVN+UastdtdMl8V/dV+C1VZjh/BidsPwgHdRW097fFy6CsNqfZCjJvLZPiSaK4MLM
dL1jxxrNVsiQoTbQUrSN30z7fqrVDPPAGrinNnz33j3nPjD1rwIWi87mRakmvJZKOdVgiyT2wEMU
AuZLOmhaNU74bsSoxiO7G5T8+2/8VTeACxGlV6SwQzStP58XpSP0Kpf4AsoQBF8B5mC/XEWNptAF
dLa5EIDIq32NNRErDhnPAFEZBkqnABoEWp3YEUFQ5gYH33AFyFp94qcm6A1A+26DQOOF5VZVXJ7b
YaZEaBzG03OTQpJh9xyv5D3YSsRxj2pfY+McbDRHjhBavUhuNgBIMV+h5U8ueXp25CHUwqTUYYnU
1sKC1T1gouC4XpBukA8sKX430NyFp4MArcUVXtbsR3bp4DuCULV7hDNP89IgjRuDxjFet2YP0hQk
xDQio0rdt5VSLjpcz7y7w2CUW7wpqTdE4iVIr5i2KN/1UNNaOlmxz6KRejd+OiZCB+22Vh8wc56d
8Ha2hI5i/cs68luefvTX0tU6fTzAiF6BZL8Y0aBU7MT0ZETSI6IbJR+nqUbUOx+E9BJwdpqxOKXY
30og3d5aHGQTMEyUXYgTU5USyGqdKLmkEW0pYODBdLKrWv2MZNX+S7tvDweyxXypJ0ketLNfLl12
jEXqQH4tTMs/40jGQJVSl9A3xkL5NWT+Rv2GjyXkXSg983td/1oBMzUrZhpY5aQf2537U/Vjou/X
wIWcraK0seq/oWc+y8DobBXERjacznbsaDFekUYX4EAxMR5V8JLfIiyubQPrvBU3JVtwN++Jnh4a
K6bHEShcvWER4axSwhiWoczoKxnqf6M4Fk0ZH+TFWSyFLyxeOFuZNJQJTJxpj7lKpl+wNDCX02ls
B6KNrYxQiqc820nJMIELZ+U0H5VpC7LL1xBIK/QcM3NP5X8UdVQyhEVOHOq59ExZ+wWz9RViE5c0
Q5ifNn1leZxALK54pD7lpvKeE4zyuJKLf9mnzAUQ3Z/CQ71cm6WX6GT2HsOeLF4S99s=
`protect end_protected
