��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��)�/iA֋���E��/CO�H���O*�#q52	�"L�+��:{�S;�-'+���UG���?��>�q�:>�}�8%V� E�Y��Y ��>nOr�����fO	�v��D �7����')眎Z4�!9�b#�5\a�� �l�I�a~�[�l�'��*�>��.��������h�?��r:-���$ٺ� Qh F����~5��K���6c��� Z�y�?g��;��j#���)h�k>��ڲ��X!��pT?Q������yf܊Yis¼����ُ��	���G�ʛ�l;�g� J�ϳ"������/�Z*��+��]P	z��>YK([P�͊�{�_1#NX1T��Wd6���\�;�7����]��n���4ȡ)��Td<ӔES�o���!J��G�Rj�&� �9�\��q¡���%�稼Uq1Z�'���7�7![b��e��)ss����|�z�� 5��?�UCou�ֿ�*r���b76����1^����[�Hr�:v<�����M���8�EmK����:m�?��O��8�&�	$qf��Έ��i[�7o.�U���ٰ��wA�{[��Ah8Ƴ֪�K0^�dϒmL/�P01�o"=�5��Pq�&��d'���}58�t�W��ڔ�/+�q��I��3�����$� N��f�`=)M!�^C��F��4_�7m?PQh ?��?Q|d��;��wn��Le��:��~E#x�d}0o�e�|���p�37�����)j��o�N���bՓ'e��A���/�]�:55ɢcp^�{#��L>�Y��H9-C���}v���7�#>[�`T�^���y{GmGoA�7��8;W�o'�/h3�P�+�WE�n^KC%˪q}�T����/*�CN����36+�<��U<�<��!��N�Y����Ǧ�V_�۷����Q��L���UDH7�M�h���μ��o����qe�k�$q��P�G��%��j7�Pr�z`T�6OB�?�M(L*Tp	c ��Gg��/A��/x#*��}R�����$ltJ7w��X�O��;yy���O��1�y}_m�T6�_gs=���Bwx՛��ݡ���v���ݭ\�u���r���Fwq��g�TM(��c���<AQUڷ�i���=0�йH(�@7u�2b~��J�"�V�(�dȘE�l6�^��T���Y3(.�"G���u�'�˰��f��1G)v�QZI��U��:�l�^\��Y��Nt0�ca90���M��Q�5T�ϐ�q��b�$�<�c��C����G=�>GVZ�@$�+��HC�q>ܳ|�^B/�r6G
�Z4Ƅѣ���N��$<U�*�T(�m�5Gf�ɓ�v�m7�b�鹷��z#%�JM{�F�,�ń��xEu���	/�c�rz��TT�Z_jh��׃RT���tЪ��m�����n����%�=R;p�@����-�;��	�ЇK/я6�]�E�	��W�
�g
��1�BH�@r�ݷ��2��˶j�<��+��+���kЃ�(Z�b��4�!fXܶ�W��	YD�S��ϒ�Ou+)���s�Tj�?�b��\����Em��mIY��t�ˢ�D}��|hQ[��y�lu�U>��{�H����~rZfX�ܳ|	�ǖ�C�rǿ�@K'��Ű�f�6�re�,a�,�Џ�_�/?9g���+�>]e����кȞm3��afqT3��[�g^�9�ؠ_@.F)Hgu���t1z3^X�y�yО��:�!}ޝo"���Ċ�y���t��z?�F3���"����$�J�{�q���Q�Y艋����L t�C�I�Z�=F��������1j<$o'��\P&p
pq[c�X� `pr6�������y���%[��b����Ϲ������z�spY�Л+P ��ɲ�J�uc ˴K��Kc�"�1L#�usic�p���_R�K<o�5�'��8<�v!������YB��w+u&@j��u�R0�o�*� ݶ.�s_��ޭ�?gg��*I~��\���Y�}����!N��#	Y�ܨg�mh��������
i-.!(�y�����}n�=*���a �Ӭb?$x,:D��c�U��0���S'K2ojTE���(�|����q��x(��T}��#�>'5�L^Ϊ�2�cߚ-�i�v7I�%����aC���BC��R��gq�
IK�7)� 8��Lt��S^�����;���2e��ot�~��]��rVr��q,N��>[�L���F����|�ď��ai�0�ԝf*�9I�80��G����,���j� o2;.�T�0�k�#�҂��h��o�Mc�6�7��w64�`7�X9��A&�D��~��S�i��RT�`����u>p���VT���IGh�%��n�;�V��o�۳q("x�4�с2���De��>����B:����cߤ�6��{��z�h���N��\��4�˳A�^�?ZmF6��<��B,J���$Nߞ�����8��Ӳ�$�Z5
��b��p�z� qPQ��@�o=4�ϼ�@LW�"1:�T2�=��}�2L�l�Q�'4��h�h�������d�΍��Iч��������\��`��<*z0(�E�u��߯7��J�f����!�sz����H�N�Z8pE�Wż������dM�?�h{���Q��
�2� E������+V��O����\�h�]b��ٞ�HEs�M�I�_,�>I��:�5k $��5r|eC�6���T�Q&�:��$��G�dO��nU��X�N 0p�K���V�����HI�{~���[]����Q�DM}t:��	8�n�xhY��"v+�q@5>��9&��QBޚ�Q<��X���y����e^y�ylrF �P�MG�1���B�c`P�`��ɝT�K�%$����Cf�&�+��ګY���}�v���H��/wn=u|�iM���y�fۭ밨L���/��=3h�������w���,�뒾�>H��=R��y+�o��jݲjC0��{������KU��Zᴌ3/]L�Aa�us�_�f���P����`&F٪��u�8x�0��l�@���t��o��@��E��M�5s����C�M���7VK��?]M�l'��9��I�����S�d��ȯ4}�|\I�
��sb���6o.���mfz[L�1�>�&%���x>BG�Nqc��g���HK?�&�\��T�RhG,��{�~�"Ft��\q��<B��FV�*W"�J@sU����r݁8.�7�Rh;��+���DN���f��]$/�����ܕ�g0%s�go���wlZ��W^�1�i+�����%�dM,�F��J]�݈x���E�s�*䇧j	k�F[��3]N����\�ӹ6��:�ގ�i���|�M�>�Dku�Ng�Zz:�G�S[ѓu���lp�)��;�8!��l� q�F,����ٲ��#Km<n9H�)ENޚ�����>�������4`�51ʫ37�<���,�I�,m9��(-��[rU����&��M�Gw�(5I�B�,���1q�Fdf���S?|(�7S�h��,~��=��c/����',M���Lzy�ky�*���!�>�
"JZMַbG^��Ceߐ�G�!��R�CD�����Q]�q�l���9MA/ß�t�9�{�1"a1�2�k��$��櫴֡NW���}���P�(�Eo~�6B�Lo�uk86ᯉ0In<�E�Ja<��v3I&�t�C�t��3.Rp�J�<W�R��9���X���K��(M:?\��]{���f05O�
�Gm��YG`���M9(}��qL��Y=;����/).��?�V;�`�	�����uV�����������o[T7��%c��2"pxd��X����3���t��X"�zLk���ο6�0��κl�E e��'�{�^�F�4��r���_{��R?���o��S8)"������� �mLt�Q�%�$�N�d7�s�?O �>4�	�I(�SƮ��*�e͓�Dw�S�z�Z0��w]���rr��q�a0]�u�*�a��1\-�{��+tQ)����������	�}7i�L����;��F��œX�0�v��A����{a�/�ɎW�����d��Pł��M[�A��!N��G��A����W���s����2tȠ*��B�+�8�]��i�Z�Й�	
�e��r��ԕ����.4S��#-�"�����湤�)�~�}�_`��[�KU� �_eŕ����_���(�����ɼ�Hw-�� �+�h�e[�0(�̻�f�"T�	���z�:�X�HSa��'s���ZPc����b}��������P��"���T�/n���01H������
ǖ��z�A��ͮw2q@��(�&U��X�m��>X�j��G	��$+O�\�/2�����|�����EH�e����^WW"ӢkxT�m.\-K�q_��1�=�[���g�;�1P%�Z3�H	�"%8cԓ�t�\ ���CBW