-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FO9PoDKYktSFEHyNaw3dY0qArmLzXceQFvvDpF2wvfPlRoM1+8w3HCoQglJJ6nc/l1TC6a+z469u
6xsm7t/MZgNg3nvE5S0Gs8mdHDCSyJpXrQ0l48BnA4geYKiXyMhVRkB9cZFpn+Na+wj/A1/HRu/h
hS/q8pZ7rx/xvD45RutOx6b8BBoS8bKXz3twgXcrz/anc6bKcPU1DHQifKHf0Z1G6h3W/Jfauam1
ifGDf1Bl0P/i+wcxgdvbOhMHLwNg34b93jsJNsjrjL+HqOR/fuxuyK0dnTXf2WdrXCZDl7/yfH6L
yNBVpjdTXbUYpI0ReZ34VNnjxGhFhy8CDyHTjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8128)
`protect data_block
++L1PzPKUfn2C1GY1xT6SPlXLTWypaquknrkH/UoE6EDUvqxmVszWvXZwp9aZDfbZClckdfzyW2I
qp+1w0I4hZdPkvwPYE+NoZ/gdVEq2oq0Bj2trg9FuuBHBNdeOjYItyrkFbn8/5h8wKwh1bZCFwb4
RQ67VUWFNeB6JoOKljhd4iQY0pF0JagdMcBipeJsBmd+lQKXqzIDFRSFNiGXE6m2sAvmBPMLrxDM
UPdXa86F9IS7A1VvIAMW7mcj4vQ1RkrSKHbcF6BLj3IQ2vTK4xQNESbIug18EnZPRNj+VjW3iogp
IWN9e0leBhqpIS+yxsyZHFUHgJwCvJDyZdAqTMd2UPBK3lJEa9zlRe+Cw4+lXElU4M1mZK843uMg
RJLfPcPeXZRL3leVdt+4qs/lV3Oen/sewmRxaMTuq7vFV7M96FCoKylSvscno1K+0XGRS5YgUpcO
SmJZZZljTXUU2tH5qfqajBXUmCDizeKD7EAAApUZ7brj2KO3ThHE1At4eDOE2cFu7lyareO8yucM
XIIvU4O6+TxDnha3GWLwWIPMxUMXztku3NTKaDcyh8ugZaWIE8PCryaz/NbGsxmEbMUHWfy4tIyf
yUz/VmCGDLT2DpOVrLPgirz/M1RQTJsxroi4xN/4TRPljeML7eovWHPS9V6EICGu8o3Wrin+M67n
03XCBtjyzbuRVS59VbYM/XpRLNfoQlcOHsWj/x7PLwV0gyQHx3+w0Z90KZYbQJnAwh61Gb1XiMmO
jTid9ui4ZIYi0SO2AP4Kkw1zd9pNT10zP+9Lr62OKXwCnIPOJYJ5pBGiU95qEu20Df90ca4fNs3R
c9jbLcDkVhEv737EJamIyckE+mKjGwI73fkMg/eYDqeoB/9c8+yXbFF9d6318DHmd2nBKB/Vj9jr
gvHE5VGAman++AfyGfm5yD1BNWWP8sxghB2vS57/bsJd0jrCbnYvSlWyxn7fUkv2CXYNIW9OXamB
m7oxbJOp/+eegvAdz9QX5WpZNYPS34fc96iKGgfNMu9bVycYDBz3m1SFduBh2528yAFTjjFAnC4j
GAdxcfl36Pimi4eeOLWCPDXgRY3hoOqd2RxlAajKY/jFr26vhoBuYpxChmzYrnllvmvcym1rVqq/
9y0CCF6qkuXq1tS5OvhM+o+UN38r0f+OZEMlS0XPzmUYevWaIaf6gJWvm9ZYnNkbmnyadqTKRsl4
cY5CN5A12CryNadop55/guYgcu+R6mjgovSM6X6Bq6oGNrK5Hz3A6zJUutQrIF1bD5Oz5JAm1aF4
oAR333uZfHXman91G8lxv2Mq6dAJCoietTSqMtxFR4nbY4lOpuTRFuwvKcwM36gkDYqcflli8piM
aOZoY3UBm56FLF9MadWB19iaimqmecsGahy7speAUSG9UeWdxJQ7RjOZN20GxqdarBDJQBO3JLvr
Ylog4sZOBGZ4KrpcCMHhU3VmG698QlapdeVPa3VuYmaDoMYOCJwqGM8pXamTS9oKpAQVOkFhhhuI
O9PxPQYETwgagYrkU8/WJNq28ty+gJZw0DOIum6yXA9X5eYrgCR19WcsT2dDYzGcmXvjj/oDxBK4
Ws+kmIj+UsywcZL+0wnYv02XYJ7ODeF+NoMSdr6eUfNQRsiwt3qwvZqBS0pl+Mb8fEOtvVnmjZw3
vbq9IKlJQxQdcIxxSElW0lsOVil4snKTZ2LXsH1rd2WTqse9llZdKhpLlH1hiA8K3yXTlGyMZQ1O
QrufMNavRFJ4z+ap41o7al8E02iB3KC75QHUAP0GOHSLe07lE8W3psMnnsITpeg1TCCBrj5WMjAP
xz85ZW6055mylmP3vBzQl9MAwkEcVFDabu4xg1uGOg/Fnhy9H99kDeYaj9skzjosCblI5s1xMiY7
gJJJLO22sEC4LT/6V5g3C7efIUzvqTJBQ4hs5JjZHdy9pqBoyx7kP7awahANZzEEMRRBRuFmjJz5
QvycIZ80ZybbvtR66XlUayhx9a8k6FG9kFenSgkXq2aK6U2YCw3DikWNWv3xl9uSPr+4ayKtnWbb
PTFveftqRyTv4FZamG4z1FV3tZ/xi5hvwiPerzssGthEga9X0wVBunRnyfW8mYALN64wCG589oMz
reeZJ2uy/SmwQJDn09eMBxb4xoX+LVsJPsY9hHDswRwPRT8Yefo6Q7e/orLbA9cetS4oTmKp7uS9
VhnISGZ9ABbkTqmEBHihlme+Zr+SNiUZJs5Rg6h/3FtaH9o0cYlxlmBr+RT1lPQtqKOGjRO5GwIB
xcfWXbiL7g8ROHoxSQOOy1mj3D1zsEFe4Bi42UlOeawNJRmgGW+zESnWkh5vg2sehSbaVH2q2+aU
u/ABDxnvu4OgzBUbPUNXIUXjJyLeuHt08pxq5Z+Zmt9Dydy79UuiWhDkbuUzEA+L8sz246dkStqQ
Ri5Pb0VIw84cRWwAxoWarlqRQqft6Wo65R/3XRMAAOPlDwDHNptAZWV8rDBlayO9JxZdBh1uI8jI
g1zm05P32Hip/csdJdvJaQh7C793kWUqF70uSxAGNp7vTJqSAtQ8siAAiyh9rujEsNT84rB/MY69
9/c5ePrhzJSWQA0vgkkjFXI1PdoeQwUJtmxXn4CyHO02aoA/23KG9rouUr74B0qArJVGUsN0iC+L
S9Pd5lQAYDlbVWx7/PWKgjqKpZMaijISBX/9ky3hp7TJabeN8UUb63lZK29QUffnt0XA0a/HxyQj
eaH0SX3KwT+K+ix9+2aIrEsWeJMaugSp7dCoJoK2TntN8CWSM5WP3H99t9KLM7qSteswEYKEC0e9
NwO8uie1WV2sJFQeSAkxH51ozQ7l9BJnoJvzO+PQJ63QA9+3w2naBLItDNSwGem+XFz75Ibt+Cvq
+6sa8T6G7oV+TkdzqqIEBk7o9IrjFgFCZS8ACwWL4QhInE0WBpkz/n71zaOBj/wZcefbbqQgiw8R
Tz0MNf0z7BAxTbx6WuIX37tddwohS+iouQDawxp2z1/uXpfzF8G2hHjPgmGsE/jwlz5Id1Nj541a
lk86RqtwkbKnNiUMZnkd/vf5wvQIA+8vLItbpmIMRpRI9RXEiXYqd7Ho93wFSuOXs13OKNvF/RbK
uR4/NQsLKrvgLc+cCf1YcNysiRNaUt0T6DNVlOPRXmgUNwAEmF1j9+B/Fchpr99xEJLWO2Eu8BvE
t5rh8DjCmZ+U7w91k51J6GaoeYlt1fbds138ecyOa8bBbI1IbQMBCOBU51+l0QdEaS/xM3/J908Y
R8EYkenKSH1ajKnMkUgiLG7Q2E41MG4/RInz0HxXqgU6FaW0qcjURpzoqrTeZsbXxM34SVXVaaBg
bho8dBN6CHvDG2l2AoIeSvaQrroK2AeVxg3BI0jYemsTuwNd6oQDve9MHTh2zHbAN75dQ8eEA9J6
nm0r3o9yJpqzYIjVnmGwZaR1jIFsd8Ks6yFX6ROogYf7J1gLrBcO1Q0w7d/zi0XVqRS4WjKQdfFt
7dWT9h40TOzV+bbzI1pfD1rCUGJX0lLlTSBwE4CH9AGtHrLkF49dJWvRNqCaSKI4sasgcLxSfMGC
3NmJrR5txcllXOranEbudLAaQpIYXckOky0KX6gHx3QmCphYR675Uf28t6ILnWk0HUSxLdQUYU3v
JoRqVH8pJqeRfSkXMFscLEPpJXiAhF3iIjZtdIwyKU05iz90WJB7PgPVtVSZ+Nvi+pRjnQ7VN9/u
FBWGq/ltSTKTyssFyJu0pp5D3zSfwwgcP23yll/Sf7Hx8x42CCSYRIjAr14bK98EJJVl7yHW7fey
hTofJuM/ViDQnu63mUGw9HqMKLgOCjmTHWgO9NE7gqVnPDf+c/Dt8PkOS+htlDjY/uETJPhxfd22
4KmAnuAC8BvcHzgOVt+mC349BsOCOY1NT+TOtvi+1AcLI4lpRAw+NgslpA2x55YWoP/iaK77NTpc
065TwWTQc+dJ2AYAn7i3FB/Knhgxz7bOFQkTEyQczgU/Mws20ys4fMfG5HX0ZkqY/6rry131Sd+d
9sc0jhDZ/5tWn7mPZ0NTDbJ1Wp+sRl/RPe9kv/my0Fu7DzJ2MXYTrmNCSGNCOGB84o8/rR29huS4
7bupbi4oGHHcL9fDdnDQn3/QoNI2BGSJBlQF7e3v0J9mcLq/VyuOCl99fgGrKpO2nRjk32Jz6sxU
JT3VuGzXuksg0ea/NvFPlWtikhGQckaWrx9KiUcCN5G+ed9+S4nDbJi2omJFCci6JmusZyuQQk0k
jaSCwrgZNVRaBamU3K0YUJlzQOOHdcptkW0yarqlWdc4W/Y0N3LUZ8ADTT4LUKVo7aiSHy9FBAB3
sorpzhr20eCVZnGNGhfF2Qgiueqz1S6M0glyZSQXxcOm19/3JGf1iXVOB1ntG+Go9q/pi/zRh4bW
HLjcHcitTK1BfMzO8jR78c4C6kuTQCPYa1uSzoGLsJTY9ERSAMsl1zcwqox2LEhlHvrFKmcGPJ/u
usdyW8N781u+YkwEKBiyJiebuhnCF7iVzEnPHySMoUjQaLz5O0KWzjm/m80SIFSwk3eRdBUbItjH
Uqv2e7ULidbBmFspJWAtQUCP+7AWTuPHnS5cPMT4lV+M3j1Jr798G2qdhv3oLXUpVv/gD3ax9Ole
3IX0CLmdBc7pEAbhVk9IMD7/Lp+Uzsyd1At8XwhiiKK4I6Hrb9REQF5D/GkoRegzVMd4D3WQPNQn
bbvg26pCZvkqtEP2doyNRnEHE9D4AX87Rsz4zklC585nCzmXNZo3cBYN+j1a1oZujUgZNNKx77O/
+Ow1rxH5J7804yHcAxwvvybGdhBIzo0I4DeLbBm/1bGi3hfn2ePpdHl7XLyPRiRLfRUbgroQ1sEe
bhx3g8z1fz5mWiqTfjDNrMkBQI15XNF4wscIrK/iuTH9MgynElg7qE3/CFBKZxdOO7G77i5fSZDv
H/rahjH0vJxQMAIUamBvT6LyFwbWgTVPzzLdnbVg/2fDGxVdzNIjOuGCPYnzQslbpBuDW0EG6401
PZj+aMWJiVrb1+gALzNnDoTIwQCrmxSCPkx3GvT3EdUbSuww7730CYmTqGbJ/aI6XMUHaFZjBBpD
TjV0X1+Nubn6VwygX2gGHOXIXSSI4qiNql40aq/IABF5VWrHG74R50HgWCWX9Pmc5XOaCG5++78G
mc4exyFUJgic2CbYTiVAExrp7PkHyRxBNIaFf5jJm0cnDE7w9v90YNPU0mGkEnreMigRFEAFgeNY
rcQTOjzwIxeObOohoy5j/rahj+j+rfkoi+JeSc2R8NcCjOEoS6LbKgYITs1K5NvGzN7M20LHRNsR
N2lKcRR1Wa9f3KqARmMQQwiv3VPjcpIAOjTBvrkzHutlgZwC3YfJQg3tP6XryKIMMXogRNbjKLPp
GPvZgeAMTvqJM5SHoQwLA4b0HqDFq6r7YNupEgpyzx4IxW7tp9lWYNou8weVJcfc3W42dZtMsRqL
yXKt2cfPexRWxrheB8YOnbiL8e8UZ71grRb8890qUGWI2fUpYWLR5Q+WBEPH7rfZgvclz4PkDa3W
vgMkLCZ14vPezSospd9GDb7tbov+tigDI2UTdP/M9Nrfbton6ennfiAbAgAEhcNn2P6FqPaBs8hx
vIy2+2+lslUK5U7V5clLEG4gyuIlICc5fb/HNKf7V/Tv3HpfroeLf3fUBL+aboCSwlGNKG2gBp+n
2jlnsWaPoPo5aYoIUVqLcuQsFZAzYMl7XMhyD8ygCzUPJxBF3WU6ulr3v6r3KaBN31KhY3oZTyt9
kpj4YkLhjzF9cYY/FjVYniKmtXxxOiRUcnSx6IkBhXJK9iSO8Z3futOfcdO+745Oz71CACSry1qp
mC2sy212SixI3gBwTX+k4jyonpTtWy4LLTKKojKp5pLp3CS+RCbynBxDOP5Z8KF1IoCP3itOsoU9
T5WvtLiQBEmERCA/0LgV4wKF9qiuGJYAPOR6kr/5n30A4uKCFnsQqFiScfCIXwT8ez9dx/VtTn7m
ctL+8HvvppZhgnhvYHqkJlnZ9NTV8wwwGfR9RfBxZl7qdBnWGWT+xPYcykdj6FlXudFhpYDQTc9x
iS6YS6FuYM2yscICUUeleRuQhV5I17KbyW4rUiPTKFEFv9OnxUPLUovoFltVaDHs2Wv1d4lugEUK
uvr74rME/itxGXcGglMhBIKGHkM6UM+WkM7Rl21NfCa8oQsxF8O7Gzyg09n4tMmbnYrCATIIYVLK
YWHYi78cG6abjPtOBpvue8yWSFE9dyj3Z4+iTNOD+H5FgGsB2ul2POkvMaCyfdMc3aYYrrhPWjVn
edDvv4dAXwgUrpaiH093/dh3olS8G29Y44KvNXzG509GB2QWLAgbbge6VZN8awLJuBaSKtXY5Brs
7gbSpPQImtY8ynDIiQhDtHbAfCI41Ms20Dk/473mfaMjHHGAqgyii8qo4oO7sOlSgwBfx3rhHlB+
F43BeLF/i+D2iKx/+CGc2OUaHJ9Xn4QueNlOB467DjO7C4QWfZpGnUJfT/Oco8+J2bBuVLc9+W1e
V1PTDXP5u1i16qMbf5MEUmPLrXWIqdQD5xDtJpv+R0sxHfg0M4giBpCu1nscoyWXFbQoIEPjUpcj
gEwC9iKI4v9penw7eaHt6q7eY2+3tGtLRYCfv4psvOdnr+ds+Ab5qh04rpGKfbL6t/cBB0suBBl3
ng3smeBLBTUvRlyjiop0mls+C/9YmZ8uwJjlj7r7Y3etmG4a0TdikzLphkwVofefN2b5P44GU9b2
teofcdBJRPit6Rg0o17W2Q9oDtNhxwx06ZW1vfDt+djDauoRpAd7B5fVATMt/MGymOc6VmRIXFq5
mcsjAmpluuf7atgmxrW6eSyL7x5X0TmH8ZcNCYSob/2yUNtbK5SUp2yNYSiB4olmet84Y7/DhhqH
+ypP6uy28BJUwblMbnWT6m0xqhHu+BhL5quWOW94/MK+EPIhU2/NZrJYOQ8ELepCaL0+tzConuRJ
/ubAI+VXPW9k+QT27Xfea/+DnpjJzQQHpHeowaZZL00n79e9HiABH8ZO5dUkY0tlKxv0hT/UduuA
VBdMgGZkvCUUeAOuV4czurBuh33GotboXJZzx9TBNI6RXXnya7yu2biypM7dKy5ERJua4vkQftHb
NV8Wz/KZopbUfXepOSzlH+THsWfR7FVMPAGWSLK5RGawvEJWj1Yj/oa9HrcHi8llN4MSAH6YELkf
lXjU2M2pan/gfZ28TXR49a1viexUv6M6pz/e5oIqOx92hcUQH7bUNQx1QvJpLoGiJ2q1c0dUXbfF
7FhPvboJrWweYJjVLndRZKdJJ9URZZsrClIuiCMKwtdZDt6vr41CRY0kNu9jhAGEneSFBQ01lwpz
CKiYoVaIUmpFnDEuLrj1OrG0fGiQYS+tCEvsu3XFSWpcTKIP7WzPVCPEGyE9XBn6Q8/9F5nMn9VX
icQnvLDRaQ+QOZ6Jc3nidwn33M2kOU1oDzZhMbVBfl4NABdCsok45RxRViV4lJIVVNKr+nT8PMfv
O4CjWHIeQN/cCd5gUWvtWejiIljdrvxMcvktyL4F2pdpEAS0TFSTTfUiKnW8jvJeb6/q08zQv+G5
Kq3V4tz/yOrGyYBPPQCjnCDylBMjLOUnShXNSl6peiZANN7KPmQP8BPde/WBLXCFZiJfHc4AjNLO
I51c7ZV/mPwVB7soeq4QR2ZR8mMkYkALILv3InU/Ya0FuI4+4w/0+LSKnAHcsWd+LaziN0Th/Xvy
BQ/Nbevl8RiL5YOwIOwynYI7WVT7VYyqm113oxgzEYerlk+KcJj8RbIbct+faGJ4Dh8itsDnRLVY
LoBoAREOgT3WXd4bWxOlSCIGy4WySHYWmp/RRrMwGe1GS6HuFymaIUWHrRyxHy5+nxevOfMBuxJJ
F0JqNYMt2BFxLj8G/qlIOBo3N4BOpfOECSYGxjzidxRLdtXWUBXN8MAwxR1n6I0E+cUiIGhtKRTW
ltcbKRjvcpxucNcYwbxI+1ky4Uws5WaYC+n+cCSBvKjeGmctda6JxiBEgd5VIw957YMwvQ6jxlgZ
LuALjTtWRpW/JlcZPZ2+crHbObCf/ZnVvJj94RYMQWzY5WrozA9Oq1GWwM6zq/751ZhBzAl+ZgUi
0whVcO7IZkcbn0IsBchyXBZOCEhxDZpw7XLpLgBrynCsGgFkuUMH/2/tZhGuPguH0lPuLaA0hN78
ZJgH71MYlBJiNUFHtcAOvUfU5ucGVQGYexvCdHC7CILmInEp7wqx++GuueTb2Sute/7UNSPmTbdI
cr8FytAfUrDpK+okT9TENwoMppZ5bNC+VgvL/3Njk5CIqgJNo+RR3exiODavUyd0nR4eDBtn9Qqm
E8TtiwKuF8fMT481khwBSvd0VbD/MDl/LUjUgGY+ZbH8MnKExSJo5LkN0sanpDA1QFv315z7BmWg
W05bKkRo2w7fg7pJOLq140hZ17W+/quJHCIAB9OzGOLfzK5Yx2eJF66/OKo4NThimVPbYnWvooix
DaTCPRyErcQpg4w1l7+9pxolJJz5ZHIglscBAZUh//gpv2AFQnhnZLupLN4NIOKTrAemX5W88O6z
gaj5Afg1V3OE2pnnWy7hD8dBKbdqI/Bt8KuerAO7/WZ4g2vrG5vDG1fzPJNJ+ypevtXy2CMo/8aj
MSDjAq8kLPsRRdG93tWsr5DS+i99riX69imc8DEg/s41ch0/AN3zUAKGDp336BXERjqUuEPUkRq6
usoW/6xNmULg7e9LdQk0CKAryWK/7ncTl1R204uk2ppn5I+bjBpbunl5ebCvJbW5C92t2NH68WAC
3LkseEcNm75rTqjZ1NG4AYfLi4q2pIITvG7jrBEZeOa63PdQRbBQ76XP4vnSB9I1qbBDd0suh86x
2CB9tpan7WHygu56Mr5onjt490riPSUPeEtu4/YP87Flsw1wCoaA3zHFZSAVu13K7grt1rqlGJgE
4mxx5o3o3j7/nYlowuYTMFIfKlg4Bynsud3Xzg/wN/6BceddM2Jx8oyeT+cqJMBuvmVzjdrKUoj0
l419zD5rBRWXrN+spsRI0RIrQSKJn2HSaf2X5gV7GAMjXfhIY8/PpbFkVRBQMMgARp66YnSgEM6q
3fp1D3/g8pgnTJdHlTM5dLMGljYBCFrJw4GBP9TtOEzlnGj2tqXdsiwayXzzQl7PHdLkbJsw8nU/
E8seUGAj91tfpKtpjG1LyOhpvkOs5V88yvDM6Ab3XuA9NcU5PUvOVNgVKq7HQhKecZBaWhonsybt
MsQVQ6b2zQbzqAX8lG3gA9YEdQKTTmzE4zE808ukZ9IVXq9H4ha2k6JawC9KqnFQr89yCCIbie4N
L9qhrz1IlivoRLTcZG6iXgB0ZB1s+JfkKz7UdUwBNpU97WeY+pmfdq1v5TSZHjb4C7+xZnPAxMyj
vP1uqpSsFqzaWCGCXqClKoFbuGY3DFJ9IVZ4yLO0zn+ckBIn7gd7zpqTj07moXlNqi3odAKQOPYr
KVFUivFg8H8wV8l+yqZ5WwqUzbD35OXYQPwbbJ26ifISvdPV0tQqY4xxBGqZU2ecs7CJ9xY7kMvB
Mvw0VJhBIOAnp9iW3yRRcgJAAX8CDnL/6e9niKt8L4t5uR2ZlNpsPP7oXRexMAuSBF5NrD9ysLNv
vMTBsu0+NIFqmDMg+RdcXfz1eqJEfbx5P+DzLq1adHahB26ciJLRK/Cn8lRWpXOqmZKzs7jHJKQI
inqrsv49KVZPqhwtmBxqIYSr/83NJ5jeU2LMQxYvDQPomzlIPxMJmw7XbFuG7Vi2LZoBLaGO7C2N
6DfhEXoFvsFbdE/5uVRpmtdqlFp7bUUOnlxKearPcLRQSGLKHaxiM7MLRVgQ6eF0gdACkJrgQR+S
5jOtJ84/yDsCs4BzXBx3Zmc2BRakTQLuHZachJA4WD72JKQB1EzPFuSz3ekBws6jfy+czED4NoXx
uF0GugCKkueq+LWA9gil2xWTyvAe6uHXtyRBf1/ZAcvYO6DDZG9srC1ZTG57c/gMMB9DE3xlGtV/
KwQZbZjT4hyJ3jw2exqlYr99+09+aSAXTLaFH0lr7fR+n01YaAecuwz9GkrP7LS8UOvHrdMD8ejN
knBcPLHMmCMX9BDEdtU0HbmC8Ke07rkO8ilU4ZP1bMTYrQNE0TysXQ0skM/4rhF54mDDhklQWZId
vNC4p7lnonN+DrFfkCmSX0p42jl557dHIkKqQdnqQM5ATA9BytBd1monY6GyJFeoHBlHGMtAfQ7s
iiV7bcoAbdDFKUx0JdjVdpETWqvSSZZUtdywMdGZvdxzXT7uSZxro4KXDpli1kPZxy+vE4UIIkB7
ukz7H24daiBKY34rVHyep4RMZMFDURbvkB89aco+2+00KOmV95G7Ja9TxKSYxY1iPr6t8KhmOQiV
LBhqeh2Ulqa+0PIiTo4pDOdjd1iv7t0VOGp8BLBfauRA+tSYyKsS0igaFKLDVXtEa9mtHuy0bKdc
klPlcD7lSE4TWCk0jhpF0G7C9sqhjF1NQDFvoI9nrK23LcWbMzlRRHyKU59Gsp0Bc5mfM++VIejW
QXjqnxFICfIEPgb434XY7hs9D4m98TPOp8trB+e2CH8BZvE0CWKP/sKftqf4ms00A3Kh3chNG+SB
v3Xx+J8cdLyJfeYpMe2DnasOf87cMioNpd2m7TYhJt4gE93Nh6KJR5X6HpohP/Gzm7CC1FBf6dVG
x0/MODrsiqWqCQ6URiM88FTvlNr3TVhXwqUKgtK+/gIAbKiQgEAvoG5iEvZPspsxlQruUUqvBDxe
tK59WInhnScv/o4uvpp3mLBu6qU2PCNVqqgYuJxbP/3vYA==
`protect end_protected
