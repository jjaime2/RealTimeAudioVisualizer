-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0yDEoNUbm/sWzVovUtQWuS9Eobgr6BRjJmuJHrJ+bMd1+n9I6QA7R1hzJSO2NKjoudPJfNqRJKRi
PR97p9qcP0zQeKsgdqahce7k/DDzCghQhGhCElb3Ya2EIIRLdSc4xSjzWJYb40slkNrecamDJ/YI
T8xOLlXSXcI3/6o9j51uqPkOspMCbStLe7SfvBfBBKz+ZxgktQ/OCh3Ek0O4nCsm3Z5IsRDki/jS
l7ZM/BBACYwL5/NBh3vww0LIySaRf6FbMGQC7pNdqVeLCbV4cDIpruV5U1RCJVCh25KG9d2r1vZ/
WQzcI1AncZvq7gePryJ4K+SdNONjUqe89eUyOw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10144)
`protect data_block
U744C8q8QXXPtuDYm5gnqa5Y9tsFsir9qsfStVxdiFGDjz7kXrs1b+NjZ1OahTZSkADfqZJgg1F2
k/DHA2MxSiqbAyLipN9biCY+dLX0MpwxC2yKiSrWGhDEGz5y3yIFoX8wG7Q+LgseQn5eNWUwHYcc
LNKlJl32nBc1H2+QbAUPQwz+Az+ZDEDJAV0fyXJQm6qFDP7zVENYzIK1Ew5U6JdJEHNwoIxhtnAk
4S7RnMRSxOoZ+Cs9yLgEimN+6bEeGPhhNffjsV+P5DyOMPYu0YUi5270r8wMu+Ezfne5kU/O7kT7
3El2ZmVuz4kkERa41BTNYQKIIEb3Nx2kZVhZtJByP1+1gaRnAsg3nMgFI5ASyNozWfzJ8cZhNEY8
q650ia+oUyEiN0Y1MKrCSqi8hPl+OK/31iuYTNyHlWHsLZuADKAqmgMWklmvUejFwulPYfEj1NZM
LeAXSY200cj5VE52/O/1LAVNO798CVeUs+kY6R/0CvAuOf+4WMtntk6YqvIocI8L2yf508CFSUQj
jii31GWiY+0AEPNXbIu+6w5GjJIZLsF729UOuFYTkqKeXjmZjlOKn+n9KdM1f9bmDv2w+K5h9JJ4
0JcGyIpdb/kziSh5vsUwZxxGcOEx5ra7GkErHSG12GkgcEDLLtkcJPTj/do6ewsJXK/GAtrxuteS
7HDL0MCKOi7RZIh4APi9le60Hr+kCLOlZ9m/UFo7nJP+S3ervTIzIiP0+kvMkrytgS5j0PEwfcy/
C8G5/zYVWgGedveQTRVq91AA+SAGLCOjme1aVoAAvqgvhHy/EAlfKUMuz/kuIdUOEEwJCCKAjYH8
pUdf2L+D8NCFDMUbWn2ArMn0vanFq05FUzFs0IEUzjXpfg553m+p7OWveOBZ2H4xLRGIO03Bq8mp
5DkUgLIvhef57n5Uv4UlUzIh3SMhHNyVAmHZl1gRHh4wOGEtT/IQz90+EWjUwSFyHoZ7DN8U6HxB
sm/3xQtO82wtMSSl58xnNCXdemjn6RiaGk23qje+o1aXHD4mh0exodcroqhaKE+4g9nS9Q20+W1N
nmdtfPiLmbbbF4NL6f5K/S8rP5O7ne5SogS2RYUjQHyUPKB735C7VQGwMiAKBT528tTXHyrdyUhb
iQ9YgJ2H2MJQi1R61QUChtC6WyBNEzCF1csUefJDsZzSjerOFMeiDGdt+LOQ4jo9YXmZW6pVFS/o
GwKfRVhcD8cm4K5sqfy/6ZBFC2OC/m/GnF64/DaEmIRY8NYHISRq4MqDxA26vzFJpuy3ZvyeKPMj
PZviSZ465Pmxi29KeyZ6KUVlm8JkOrB1XvNGUhwUozq9BQxWNx+x0+6JBA55xP2119AmdOPQ2Hgf
Od/D5kcuWdFqyJphxh9xrbqCGEVadBfJYImTvDZEFbfI2tfWrwFqLNxPOBwV9iUA+ic0RT5Pcxg3
/S5qM2WD1fxzGaesJ1zBi1zzq5nGwEIZRQYZ5Z8zWJYzdeNiwfuuQemk+XDbr6yhB5ZvkUON7iK8
mOZmSPfCGhyEv12YHButsofGpvE1WRwFbrg6qh1SmA5lkRGuYvr1JO5pUt7poMH4Xj4ZoDpWO+/P
d1Y0pn1DYGP+27KlTxMsyW9c56Dt43E5qsW7JtImyhj4rxeF8e9uS3ocAzAeGvyHTbpJjSQljxoS
dm4aNpDpHa9HQ9lb3ObRftQgqTLYJpgeXa2aLXa+34ek8wKBIgNxdJAdnZbjsq2axtqD6ym5Uq5s
LeOeIHLcodLMyICoBHhEb8nDXukbtXNmv7PljP23/lbljeWYPIHh/Lk2r6cAbBayFQmk2LBFkGXt
eVFP+e3ruqUs7N1BM7KDpQPpBsIZk6BQzQynC9SLTpxASqAUNY5wyLIIQh51o4tBoPgflOF7pKUN
4ROT8Zm5CgkkafxmtjM9h/pePRTkUNbpQ8Y4wYY8XjzYc5uF43ghNb1/gHnyK98uXyk1Z/13djif
fV0Js5lIppXk2qfwoGc1AFpvYSEfclndBa+av5N4H7n9X0QwQ2t4hnMBXPtVZTGKjId0wXasQt7P
NWmMfUJ4yJtrUDAIb1Pxy45JZASpXhrOrKlfoE9Bc8vF7pEflk8UCP1NWejCipxMjtpju2F1wRcT
x1n/cJMdKGW3DT6fz/N45jm58av7peeQPfUeRzBl7yzTDm7AAQFSVSY31LP9aeDYhFzlWU2mjynG
e4s06vVNRLskrgZ/uxy2imRF1I0lZWB7HnN5tFPElWLC4urKUvFrsijh3V868CpkAi13K4dvEBxt
FaJTu7+qrp75Hpp/8Trq8MVBu8kNGUhCyxKi2PzU5q712Wae2PqoV9epqRpnSaH9SXDBIN8sYSQe
a23wWNdDxeJDupkItJj4mDERdHWck6sMt6LlH4UKV5g1DO8xWQ6n2kFPZyfzfOhcuEF7NO7FFV15
V0NWtLfAwwrLS1T6/W4Dbb5+oGhWjJumAO+KYFT5C9ZRu0D77D6h6aBNc4/4RuRGuWlKpyyzeKP4
fd8BqvqcycOE8o1hGud5ltnFBqiFJTacTPXFqthK5wIsMDc8CjwPMANj1U73PmXgD7rnB7tro/vZ
A2e1RFQTLJwqfehfq9ArD9FMjZRnUCm4E9mmZquHVH7Jm5jjlT/w6S1aufC7ctxVbyxtamlhYDPP
LrVOFxW6QP2Wdlb/XvViSD9TYHZdLeWcaNoEAq+haXkDtrm5AqVof9myJ6iuGaxX12eRCyMY6luc
p70R/3GsMsXAjDw9K6nZRAP/fTlymQf0PH3/8TiM1U/MCd6/6iLv8J7nlbh3LW40n4h+2/BPFoTc
9J/JblxG/LhO9ndvES830X3t7X/Gj8rGjECfwAoM+fKtPUlK62s1V8USH9l3U+Jd/h5ZFEjrZQrc
6q7WM/AQ3kLj1S/SKHbDF8xvGH4YyOde56bgvBQ1oRvDl5eUo8475U6ZgRxHxh/yNOobUzS9AHOM
DusIz4h9DM982QlU8wSBm4ap/mDdnn60Bn3cDtHsanfFicDxuljcKyblc8oek/eTx3DD0oapvecW
cU+/VsV60+5yNDYTqTTJGqKywsXQsSVb6E9OarJ424WgwZuktLExy/+wCvK69f2WsP9U4PEVceCm
sSFeFK5/Af1cnqH4Eda6hioSkFScdHfRhANGJ5OqB08ZU1Blub4iI6O+2zir0WfIGySu3dUFjZDW
a/u+tyfiiQVYWSovX2FNgVAA6rxxIW8qjOWsrNOPZ0CiFPe8eQPrEulFTFdzzUQEdPG2xrZiZaqx
fomU0vJnJ7B3Y5EeCLtPsSrMPU1ALQw6OTX91HejmwbcG4tFCSmOjWIS7y8SSY1ZrIfE3fUzFZvp
veOfRkom/+zjISyKfJCSPg6Jkk05hrI/mvMq8BbSmmXy07PBfbWIdCJ6R7Tq7UJRDNk1gggfrIz4
m1Yyth6ndcWDc48hi9/tjjb+nh7Zt+b/BqZVdZKx2l2sjVVIDfa+RzoHq6oUV/ox47TCuTYJrAqE
Kub7tBsRqxQxGhYqBaF4NVBBPNmD8SXmW2eZtwmUgqSeqd3NxwcW0kg+ax5WD6WoscMsz8Zg7Rq6
046CgTrDaF98zDosHkgJY8Jv9AeAYYGD4tugQUr9/VyAVrPp1ISsO/WtLLraxdd3lH6w5yGck7AF
ZfT8wJR7vsUu6vhQxDnx/w6m89+MPHJg1tInGpWi3IceISSA/yg3gMT9wnJgAhBW1ngHnlVov8IZ
5KBfVSdHHDnAx6DitCmUt10SyjjiQje812HkixGTS3b0Z/tkD/Kle0Pu3A0mhzd2yNJWa63yWYeM
+fjf4S9Y9PLSTnt9s0TSlZWHMq4XbsJOTM0cFPofZYBmjPggpj3vgdsBKNvjqOsdYdGmCQL1zrvH
ICiZVq9VhuXOKeQkWqypxo8D/XZ46WTGKC6VoP1vWB8oj+BjdeIvDYBk0GyJEbnqS8mYBt6NhDIz
Kk8VHOpNGOJL+xC4XvDdSbG8ILP37M/tnn1w7mENuMUw/7pgn15iA3kd9I1yMCKkQ9R36WLoJDmq
RLoCvQtdovvDjNCOKDOieYiDYmr3RFUUV/y92QZDQ7CTFdOpG78FXznMN8f/l7mVehES9jbRKbU2
FUz9KcIsLV1N3ocuA5CobWkTtO0aZquDYdoWtIcopZl/0Hp2HqRpWIeKhihGuj6H+05jIIXbZMJH
pVN7ieBaXReegU66OjT92FhvE+owwNsq/r6ygmwVcXEOkomCnQ6JJc0u/sGu/qBx0U9taTDKtK1j
e4c0PyBV73yogBMVFh3zU1mTeI3rsZUu9WKuVWtHpkxMSgMrPPlKsGYEKlzLxA0kUYMcjgafjlJP
D30DnYNabbhpE1OJo8lrWULSd3CrgqWm7oWp5ps/0Me1s/SBu4rdhARQ2LubIOKo15CYtibYVTLX
Myo6Qxn4eN8aHX7r/javzCq6F61CKb5Z1RpN5rR2TLiPsnX1gi0GK5iYnSJt+fnGPeOjUPsXUkTi
2zXSSdqxXHvoxI11/IOeO04kdq+qcBamd41UL4f4SvkdhyJ35own7VU9Rgx9AzQFVtBeg01gne6a
CMQcKCSCY14DHBMgGmiiHS5ifqCE6o5He+xdH/TVcYmhXtXvgGaoiT+MCS6P+VVJQzz7AejProic
GoLOx+bxGEkCxQT5DC5tZo7xSQT5clZIt084NYuU+CDgxwloj+G165J5Ivba3twcO0FrpTgQL2/r
YMxvQl489sPaHWCBCVermFpQkiJbfEem9je6YXJsdr1rYhobYwDFaNkQocQRCKMs0YgMOGLGwP7W
4JuYAmTZ+B29tZb7qR9rFM82tq4EdaQmH7cHA//tATfB+2WvVPAYjghA3+kkjXhGnzeuBuYK2sRU
BnYMjT0EOqEVbRsmfZwDddt/ftO1xRtA1im3jxNNkjg1f3e2+srEJHkGgdE7dovjQx1XElXXZ/Ay
JSPmx4E8n/y6l1RamdJlRhwAOnzf4GYMxey8/1DV7nHaFJTjxv49S554Q6PB/L7eZUA0ZEmhb3sX
APjYODFkclzkm6fVVlykiVAO1bcQeEP1MgxmxtHCmcssro7aQBh79780rgAGMvPG3HB/Z9uc/ykN
Vc7HiDMa8WAGtJYXMdEkAjSoP5nL/FVJR9ytbUhVIUU8tluByI+GKkccYSZjJOr9xGVCWTpbIsiF
dba00kz26pK9g/3gcEevI3+BYoRrH2Uya9ejgWmeLuw6bB70bgYpsn90ccze1XCt9r4LmHjFZwaA
i5d5KgZwOzythRY+fBQaL/C2YdBVCqpCvCPAh+OJfu9OIHoL4E4pTDDwfvXmrq3rEviIOTQ3uniY
pShpjwMlNRpUnaXpSTrTSuOcdh2yqU6A7BpT8tClIjxcRKp5dmP85Zb47pHbcdkGdJTSCe3TylB2
UNCBB5LFFUCqiLC5arg4hLpIDWhD5wGVgoHwfp/hGC2TYa9orODDDhYJZtOYAxA09XtUHgIexO7a
XkddGDJpNJNa0I2d5qJPY2USLI66z92Te2oTxpw9qv2ZyWE6/StHCHf3Az+ZVt8vEFUCZffp9Vsv
C6eFi2Ln+ugyXrtWE6M38Yqoo5VFexPMnT15dQV9IxEw5aJyPGUrvGYKuLUe9VRSyp2L3YByYhpV
dIYcSoJrpGFYCuryFsboaNh39iM1hI2APwMBPyjg2og7YXkTkw+PNJTUCuceCwlTu6cCh5Or6uA5
afhIyv6mtEvl9fMFv0zS9XUOs4DGvrkHxJ6In3dWNQBpxj0gma1YVkcN6kIAAQAvRMztK7jJNXwQ
Lg3a+cMciQ3G1rdrX7VkjOJzvCC6AKbvWlRERlgShBhB/Wvm+LwBmHeeXIjgv/YEghiVJGIHwdZm
xFQC1s+nTU1jyFtniNkRaqDEQgXMWgAy3kTPzyzC5l5JsdodDroKVWUTUX37VEsa+gaoJmQDVV/W
wdKSlwqZeCe6OqSmYwFwFFCwU7UQXMK4mK/M1Jw5pO0MI6n5E629YfTQxVzLiJ7TAWt9eqnEKAET
xu4nq/Xq+iqsphBFJfRY5nTjjNCqnGHpH9N+MaatyrvqGuMEVR18Ldq+rpb4pst8zk/8XCKBC0Rj
YuJ9+mdL6s8q9C9I2il6FB+X70icEKxPxoZTDpLhr8CllTmQgazPcC63E/XLOYsJLxPurumvzsIO
l3oLDM5mJxUTwgndONUbedoY3TsWjHFTPWjjEBqDZ13hzFeEaoxqu07gsJ6WLLGSx3+Wb3uQBMEk
tnTuqSmGrcSh+EH3ovVtrmoKFgoXJvqY7ucHZnBKDvpGnlw1jKNw1JCYNLfiD8mddUszDxzDrxew
DJQWkHkyJODQDoSjJF9+FL7zSWxwKZ2eC/wD9x8vqhz4MwX7bGyMxGE3mDst2TdtDnwPlrr/13vD
I6tj5OP98Xb69bscIgRalKpTQFmEBjalbMTm0Xsnr0m2tKIKMHJfLXxpnZBLfuPNjz2k+LaniQq3
c+m78/jeV6US8qNArp33Ej398QARAX1mwbdo+AfpC39Xfw0uG0tM7q4GZzbKhAeUIvV/UKAyuI7x
ziFuF2XS9UWvhfigkEwAY6Wzo9DIdmaRpc1weOr+63ttsEY7GAqKsoi8fCWcrl6eMHqZ28adALh2
SGVrIigzTZJBoFMkmzhqP1+wYDnrZEi6g3+77NybIu01v50xVyHkhDtWrkrnyIapIHNbLE7oRAeU
irltD79uweSr643LBcok62u/nhwEciFP/L+NT5eNkBabLUygWiRp039qXK5EHTbsE8M01eEFtoU1
YTylFw5Zd+ekk2ZgiK3hN5FnWQigzSUv2mHtBLNuWkHCtv9JrmofNsscp7QEgCr12urQhy4WiSQt
/GqZxUcTL8vkgT4Mz2cFKFx1WKzKONHvcPbhCiwT3u+7JiFidcr0oQy1jc6AlhsyvvTDeDWJdUeo
7CSpMTodXeNMTLVSaYZge59wHbNZZBci5g1lBLSBMHNPe4aRXAz4Ks+cp5XDd5AQVMWyqdFNeDeI
qyeTW/MDB2FGpAK82aY9NQbgoKJyvklJvF6piK+XGf2SXEZkIUGgjjr8IkOsSFmT9IJyaGGvn0aX
Yoyw5FCNP6YLoBbeAtvfaLt0bwTch6dyXW9EO3H5W8KbBfSsp8EqRA/RHIBuvKsSm/ym103jhReU
Ryjs3ldP22PmmSuPvEd3Q7Wdkhw3yAZblEZ5rWo+Ol8bEimOyS4xvydUPgG8cgKpNBye7//vuehE
BUyAkFjrLXmaRb+X5sbMXakLjgVTysAM7KcjAWvetFIYeekuGeTpdL1AoI4KTxDSmOnJc6KG22JO
vOYIrk29AIhIAiBfX9wHmkKanmzEvLm31CN0VfPH6QORi73OtIzyzbCzm+gaFWu5hMaRYFfFb0ZY
wIU2Up5q4rQOGWBesxCx4lXb6WNYCX6fDou34r6nfaBgOgDRE2lA237VlYwDeY7TbYCpA4LktSXz
im22uLSXftNRUIQraE7R4It+Q+3dj7K/uD9RovvYqCALeHGBWlcc+etOmipUiqKGgZa4/3Ss/6U+
g/rfBFdQqFltFC6sy2bslguxe1sKFKr1+PODNgCqThadgpOsr7Z8NUXOUiyHUoi3/0VkgiU5puty
bBKAvw+pp7leixj38yC0EmMNWIYDxtlFGFSJlIhtavG/9Cg68+c8RnG1pSNOmoI8NYaTRKYsnbRu
4Vv3ElhQ+gaJzO51nww5iIKwYriLaYrCK/XQiIvHTbDk58rxEzaPyfyapKNLZDGcOtK7uwYXMEZV
RibzQ0AfR5KhaHjMeTtgsvcYtOpWHTZ7QvreoQ6rXBOe3WKj8PLey4Ho+oOKs0WttznWCqe0BNGc
itU40q3jAvCp97IXeM+05uhZjfisi7ONR3k44E9Tnb8tMt5BvtKZL+1aPjiBMZqRSto/cxAgljdC
WkxR+x5WZDQjBHr42bI+A7hjh0SjUMX9ShWcxw/kJVRP/WTNxJ6bc52mM2T0eVDXNMIyalLG/VJv
alJMfBudKfW5fi//uSgCMFGzFGd+wPBRyvBzlo1DdQfQwoIDbjP66QU2OQ900/bwnmPjDKF6Jl+m
TieYYtcF5IvKpek7/SPD4BjFoMhcn8XR6QtrVH9Pf/fj5MIiLiDOP4321SUy7xOldHJF8ggQNxce
jMLBZZHkJ5DhFsNP1urH3rwgo+l0mHo6YJdArqLojvZMQk1hdSXnrKOcuz3XOMx13cbv+GVLsM7o
0Vd2m5eArpSvt1m4Yuj9an5wG2gZ8EjkgOmkIX+6sWaa4KmuIL0aSdAROVpdgPjubWDsK+QlwB4U
VcttY++5zfHIDlOB+QbzN+vcsgsXXisWYppvAQTsKbnnNATevGyqAdoX0+Hd4ziVm6PaHPIPnODT
Z0a6hFbperk+wcs5LxjK3mRCug5SzueOKejLN9Rseo8UZxNqXSLxmf1dq4QIXm5XeJ7xDD3/FesB
E2ws4hRIi1iIVXOAJ1OOfQZi+axbDOQyRp2PV6uI4IWrwTACLPL7YN2787eGFt79Iv1626ThOrWW
3zrAeDCaYEwivZrfKP9vyNtXi11j8YU9uE3CAk60IXPKNTBDv7FvF51Sxjlqd8RJLGoW2J93yTc2
H6EeHzS3nt4Mkw6ZUI1e/UwTlUbhBTAZkT0CBFdsyowUJVgbvWqSQCgKLDTh6fKR38xOxg6GFash
IYEHQbAJ/nZkzB2pFJpaAxqUl3TyMPqGHxkqAJnByO5B/pK5Y4/NUomFry13y4PWJNBghS5RA3A8
0bGPal28x4GLPKIPAuYRPRvtciTsiQ4QjfhsOrR3jjHe2NbL3CkUYz1hR/SlAaY8UGpqx2jTLtsi
vGRpxtflYgfRDhDgJ76jO3pYNYg+4hlhQYSIwqzbXb3ULhXAkrT1+oqIyK7uGj9hWi17+ceQBko3
/OCEbIDtrJVKeChC7CeU8ynZdfqOI5bgeg9qqxPZukNpyOgmin7v0UK6dstL+Hm6ljBKLYgIKzuc
gLv55GRXhJrGLChFkfobbO2ieWUZlkxxyIK9Li80SvV1hwEkEewtxt2yzQNt6+u60ntT5xTUngP7
EQpquXAOKFOThONOVLipiKMOQqXHZBULJPCIzs3ogsPLPD51LQFqIxBpT+rH5cGLza8/mM7F/ioF
A4svUBGm9qKBQUw2AOmwfQcx4CUdQXsqBmln7OgmGt3LaowggYlN+YZJYNQWNDoqkYIfR43gAN7k
IwI9LI4JYGx6cqfjnxxdY3sSoAH6HyxLFe28Ku1tiV4qnnobErBv25yx5vx0QXdGAxgaCooQJDIJ
5LX0RgBtdNHFmQIU/Qm1tN6MV6aUOx72HCGsSLR2U8MKIiQ6ay3UsbB+gHl8rCmIsdzCHI2O2Rbh
LvD0+cBoYS9dSXJ36505Rfdia+0RAkN3ASSsBfQQsBxVmClVfxbZnXgJWP5rjsvEggQM7idGaKsS
pnZvyy9eiEKb/4N48DbDKMjkzIYNEPC/ATv1gTbLrivQXS+wvFwdlgH9zYkL+iGEnC5JqXaPmCqQ
W03rViHHtNlD50cOM4HL1iwy2xdLpqxHFEixGhmO8WXEm0+lzXz2wiyVGmIAEpGq5XkKUG6CQ8i/
IUQbUBMjEdyYUNYfme5o9eruai3ltls4pOi5svDoTN6ps14vVp6WTwtUsBcRPopUtMjg/W4OM1kQ
PHZqupiRJuNJSE5bRXkH5EoU7drXwmng0tTQXx/D9rUfiFQMwu6d23g/Oy4kem3VB3dWvaT1SZWl
8APNtKG7KTihNrOU3dKpzVCJKJh89UasooCii07/2xHwghL99pPsWTPXWPxyvq2RIOf+uvYJogCS
mk5QkxsfAYq8JCCJRl8n3IRR29fqX7LGypcpRL8Z4ikksKziaJGFQtKYdvX2MdlXtfs5ZzSHE0rB
6kWgmYIZmomzAAYKwmWOEZ+JkcH25NME16LRnAE5aXiyYO68HQ8CrU7SrXX3ZxHUpEiXoWP/jirv
OhB8FVy+2ZrwB70xdlQUHvrpQPKvk8d9vr/dApy8Cd6rsrEgDKP8j1gPl+PudE7CXjJLyWPKvW0B
lzvfRgpofRrNS+tBquAGMum3CaaROn+qyuyBFsQs+AyFPidIOjtHVzy+PXAan4W8ZtB3FiXN0QaA
YuKWZY7L/X1cZ+JeWi7PH1ZEZD2efnORU4dJvM0mO2CNQP8P+OZRBJPf4eHc0nrcjGkHknFwbK28
yCC2pIVsG+idkddsLoZC0BOU54BP9kz+4v7TDXbNwB6/m+NQrhs3qqNHbcvEmENeRXQWlgv1A/h2
pvGSUtEY5C25ePn+ncLHu/IFrD/efit7kUb5BgkYA0d9nisV5jPQXYkRUspgB8R2W2loKHfVtzRW
vFzif5bXUFNgyLXLGqszhF/XzDt7MimKlt5nsXpOsaAL8AQXyRRpTUSvJk/dVMeyadcr5OAtISfj
CuNuWoiM3mIYUI/HWBdCM7I/0QAHpWAF1z8EWSCWqsI08vMT6lkptr2F3h6rdTjzK5Lng/MEi36Z
WD8RdzY0u9j8L+M3rdBz9i4zUellLrX0XxfqUm5StfdrEnDl3TpFKOAi12ZV8aArjoebsrJdpbAT
nkfE99fFzzXdUYamDoResELrLCD1V12sKkhjkbP0xS6Pmf1nFMAt+K0sgN6132G3q0bT4tVkjYpp
PGTxFXHZtzJKDHYkZm+dICl5aTnUWinXdWb+QBvbmqQNoPLsHPF7B8HunWTtKmjfkjIy1pn4zvu+
OqvArg7UigAoDDYav3/uYHktHwaLdO2c+Augo4n51YRGNWr5uXSaXd8rO24P1qL86VfikTtimzPo
nylobD7iBRcMEAFPCKNaov6vwNEbfOB5gd2Ttou68dTbSRhpJggyHbl+3VD9fRzVMDyueSBwIcBU
oE0te1PUrvz0h57gumNDBet2xsh4yGLbGDdX6JlAqy62embTWunG67x4FSXL7BcERVuAD0uztIFa
gp+zPIdIu1PkE/I+kwahq6kQ7xT+1yEnm/ydYX0WbftVjOq9+5pH72VaeheBdNSAmdgxhV5tJuke
V+Z8jDcYQBQquXiCNHPQlqFZe0mBpsW+SVioobNZn2c9cMxykrZMlE9KuPm4IWr945hiR7QdtOh3
iSNo7GPOoNl9Nsr8e9xeBoRSUx1yR3E2BSL37a6eYWx8gSRECaaYWYALHmlVcgNVMfHeu43OLvon
WtkIvbrkSauotLp8kLcho/1YtinNrwWiIZIzUnJbeL9EEz0KYXg8kKXjKT9ysLEGTxrofJQVUxxQ
5jy7GH0I6Ea62amEjLaIbAbV8yhVVtlFfZcch/yBr6NL0EU5tN+XrkIckoDoHUD5dhaEls/e5qKJ
+DCtR0x38l+T5gTHLiiX3RKIZ81Zxmw6IgEkJk4oiJlR13UCBMHj1QLBQh5N48sxoJe67G7a4yyg
nJjLmno6IsSrUKHRWalLmyU+JDyyLXaQOls2Z4WgAmya8gAILgEKbX2LT39cJJNA6sIsQFDdPm3z
Ue26BmNdkouF+qVtTIQtnS6LOwJGPh08uHmCE/XAFXyGM2S0GTTOQbVCF0BH2UK3/Aul5ZNBtpDT
G1wcsfQV8uK5Kia42vTjjWx9fbFhfQZnBzAXHpQ6n6OggYlDP7Rv+YwN1CWU6tJRRLYEYo7EtGS/
hzZlQvbfX/965AIWixGWIoBkB+1/o3mzRsbgd9Fp+tiZrWOthUwIDQzgvKaXNk0UZJnq0hYaSqvA
RQ6+emXLoTzVAP8kmhbNekXBakzSpjjcSIu0yOHrEDJF6dtI2peasfeGd/okUfLL7AhMgk4TFlVW
Y71Rl5go5RcCsBv2fcEHQIuaBu3DLixUeWFtyI+XkjJ6ES5MWrLBuiVIpo7SZbuvdOXURPb49+HW
Di46Dm3pztT96F0tDgOCt4XLNwUlyXmM41HYNg07ESILa2AhY0KUJOEEAqJbIFqJ0XJ8puyIIVKP
j0Xms72NS7OdTvA0JXDoA7EyzRVanuq3rN3+qOnUM43aTLuh61duSiQLZPhYFuJLoNTnjNrG8l/9
xb8Si5l+LTKyZFTaHIc7IwvkK2/kPChcasunHGFMAbUyGU43Q3yBGdrb/WBKj/100WWdb1twwkrB
Jqpj6g/uYT9kKcDYrL2GJRzJLOdlKksafIM1945QMs9MruPBTUpfOzrA5HprP8wEXcEcWXilK68E
KfAj1SUHgw5JoMtWSXeFmKDcJwO37GtNqEGpHfAzq9+8O9aeoZ01ny5zltXXT0z4r9w1paHbots+
E7nu/Gjx5IUTgv2UsABk/G3EDVbTpylPZd+9kNjxj312dX+r65dIYAC9E7pLPecTH1OWZGlqM4Uj
zQkQa/3x9ssZWhGFDSKwY+4KZEQT5YWf5OD8GURD3yVWUwv+DSbBwTmKyTnCslbRqu7iAUY4LSQ9
RlOfHvFMbwuJjnF3PWmFVFXYddy8YWokHQEJ8izvJgVJORMKEgrnRqVkEVAicDrTL318WNyF/Ewc
2j5Sp38tmdw9CqSl6/TrmoZ74hRdA9h9QxfZDqM12Y+7ZL4Ke7AdmcA0+ql6oIybboXWdyDSmWl+
6Ph9TEGSFkuAkYOIWGRl9N5Cp4JaHHe67Y2n7VqFEf9XoYYR4e5pr4wXcR12nFjCv5NrSuguePNy
wVs+5KJOwQC2RB1gbzzwLWxjlCAL8OQNfFfPTFRabL9hOUbdhr96iGvXMfQt31XZfJuswENp5nj1
dv/A+AmhyHDsiFtvJDklqXW4TPtG7km0gMc7x2WoMEh/LCvUC4J07YTxw1LIr273Kri0ltVQX5iY
FiwD5jFUOVrfMDkMEpRw9fdImVxLQWbjW0Q83DXGrnEAadfwdoKwXPAHjhcHztmZwsHpUOy7XikO
OKl7Nj/rKv/IeSziBS7/7uz+if36LYPz3HzOLtPVra9ixncXj3k33LqKuU/lcI9Efa1XdHCKd8C8
U8okAeLsKPU2YqBasXhE0iXcYiFAzaaALMpuLHYzZftS/c54Ri39pHSFYSaLIQRbPYbgQNqIF1PS
5TGKEpI3z4v8/nx0enuMkPCEys0OzZumJC5HlRftUgyIMJPtR5oQYkxtgVTqxVJTOZYT92Xl37QX
XWcrVUu0/ahwT8D2G7Q0vEcUFXMDmmm/cQJNY1OLKPgZeoQWJBdKmilmhIFDrXYGbVrH0RzUtflX
nBy/L2tGmbA4SafFIPS6te6GMJJpH4cQZxr82nTTELrRGyT4XztCCrYgYmZp/TYEk/Bk4EQvWEml
pXQiUnOad03S6xzEr1jTLEA8ftvByK4lU1y30UghLjazV3IqzyAN4ylFNSE4AiiaM/irX5/PDTTZ
R6UacF6rIaj72fzcDo0mOQdVjHsCZ8WW6yQdvnTNm9t2ixKHiENXZ26g66ydVz6NZ3Kh4ffVyR/9
7fQuTVtfY1ecG0djvC9DLVyYmUmNwr1kgfMB/CNqQCZseGkWcvmhg45SJxZXpOkriuEWc0IeSXfP
T08kOXqJTE1plfjNTqLQlADtolragtsEwSu2cTNbvPRQ2Wrub4N2NjlR4bfxxnC6AKXE1F1x9w==
`protect end_protected
