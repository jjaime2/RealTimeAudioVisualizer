-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xRwVbFHOkQRv0gc6h6Y93sYoQAx4di6tDH2VBC2vJlSgoxWs13igyvszcW90/5ul3309jokveG9I
96GIAdz85TLW5J4eYtlRvWKTfhyTluLdlpvesf4a3IGsSFUdVHCVKsRBalFQvRdJQ5tz1vRR9TYp
3DVMk8F/Zc/wDFNMahrQpBJD5xu5t0lWJvNmPbYEsF5C5NEjdJyAqmBBtrXmMxolLgF68XcGO0EF
nBd7zmtMdi0s07AwFNQnEysD30kv50cta+kJ2rvq38/zvxu0zy5tsSmePRQnhBFf5rZ3pRpDYddd
bePA2Gt6eiL1fB3VQuVaw+AfCa+zjqaDfj8SDg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5888)
`protect data_block
Dz0H4JpKjZN3aMS+ts0kJL/HAqXhRFCWAHsUn291D+zmz9aH6rEDY5wbgIH/e6B9EhvandRZVNs0
9gFqIabXebDbrOmCT8LtObLos9aYpBFMbp8DTRBxQeDrrMrh3+2o+HWSF6Ar+GsIYFAhHWSITOXH
hmMBuAej28jYILIAVktu1g3+P8/7meEKCx2vXfKH8j3uSeU9oG9Mq0EWKBgfOOjg1nRSp9pr0S8/
yuqLgjnZahvsphpLelE2OZR1IP3v5dsItRjZJtlK9/wMFzpj6/sjxRCQo1MOkdxn++XY+osSW1w1
E8mSx6Y28x9HWJ4hAlYoyX7LETKwwU9p6xMt9Hh+ALTQmzGEX/ArefLqm7fsFw2oqnEdg4E3tPwJ
OXwb8jmufdO+yks+VoznxBrY+mTruS7azEHAmJ1YhO1iEBtfIK7atvb4CgJ5VHbh5yZs9N+Jzg1z
XUhghhirR051uTSuP10fpIWz9Qv2mLQFp9aY73zy7Djyex0c5TC8HTMT5fAq9SDU725xrqdWe1jN
dUlvlvdxaKIonROoSA0li5XoDP5MCyGarQFJ8Vu4plGTVz2BgVlwK91P+MbZrArwoZeOEOi5xKDa
N1xK2YjQcRPgAz02QQB6XB4DD6ep7eBAppd1FL4tkEXhawV2t8O1N2w9me0rUn3PElgMkh7lHA2R
+P9pYQRBkjQRgDGYCH4ZU6RmPMJtM1zZzQRB6CtqLiuUHEUYtWZT5MtPJKKAizUqh8uqv1nRJeA1
JCFxkDfoNAZ619Y/EnT377YQEhVsxdktvIum37lNdwYUZ3ZvfiLZkKgLWjMa1wl6jM2V8K4aWrT7
wnNGj9kWzt5+f0nhG8NtNvbKX8rxs037faXeYcBQJeMJP6IgBgUYv4VESJdRiWs8RegGnI0ahnCU
FKBnZfw8e95yn7u8epA3iEukH2Lo/4kCSB9tcPtSaJ6a4PPSfPBxh6+XCvAoeSJhd5CwsdWJUR+q
2EAXjkYgHfMa2YglV7NLCuZgKhkuyg8fVgIK7uIcgncahTz6Fnk6Aa+DPEsuzEjNjvgjympZ3DLe
BGQSy9Nf8zWux8tnn+VM2Bd03IhKD48Kr/rWTRaq8tD8Nnw1QyLNmen6tD2LMRxldtuzCQcbOkiI
sG/NyJ/ivmrI50ZwZCy87gH/WZZLPGJAFOyTASGrO3KIKxUKfQYdz09nVT5HWLThyckNiLf4t5Uu
wJTCmc1HVV4Z4fX4q9li4/h2Nbri4A7ESzIv+VLeYXNfsqgdiPMhsocGkhYGvDbG9EmY35Uty205
KUl1bf1ChxXW0AFObuNXIvrFdmB43LgXg+pFTz/avBybS754TTZKf9t2scjeOjXdCvdeZXNsP/VW
gF64lOUiR0YOOenjxqU9v5wPcTtfrh9h+eQNQseGnEOmmjj0ZVgmXptn2vhmJptwJDX2vW8TdYka
DrC5plp4dHOFIn7mFwpM1u2wfO5blSrXCxTfDIRi6tkhCfDCwgcLaJ3gY2YPxBfw4x2tWBYGPACF
RsNkhGmIyzChXV8kIbrcEjz7DUEdDBrRrvQ7cfOoUUvwYLzBS4cMAYaPw8YgvcfTJH+CxAF33TzM
bMsfsuBV7iLxygSKrAbQN0FtksPZCEbyxAep1Y751tr1hfM8RIDZPkoGiF9TIf4tadUGI+igum/7
Wn4DD8qgkL89MoULKHAKbyQvJkgcOOxNlTbK9XuBqhaYA6e0mz7seOIKL9jHk/qFqXKaXogn5o4L
HPvmB7bSYkDAsnsKUldwaDHMAT7dhS4ZEeSAmMRqixDouXoT3T1I5UD8v936cOnyYldng/owPmKq
+xn6x3ZqDjc0jeQepNOkccqy2gkVD3i2U0GWj30ePhdb7teSfZsA2nw9JcNycqNQsvG8LyjWt69O
36nCuvUWy2AgRJMYprmVLSjHQwJLxhq4QXszFpD2Y9LTl891K77/RTPhGve+WjHSmY9wCO4/21u3
n31l8N41d1fV36oFF9Tajiy1753XXjr8jTfhMaIdLzNVFnisL34NqlIDwciPbCZnbhYybAcTm+ry
OfIqAo+1gLBWQDa1b+xM65+wLTG9l7c5UBWFeGFJMpm/WnfVKI7FtIl3+LYMeDDUc0Hkx1srUob8
PIXBZQHRhxKgzPRq08DL698/R/u9t7g0Jv+Br3WMK2m+g+jgKZsw+gSPhsGz8XX8wI+DizGwyKWc
D0dB1lrZNGUPuQd/xqDAe5aSslFAe1jPnZgE25cW6ksPIMXmMoovoCDOU3XjasQ7N/zEFr29Jp84
QpfiMVBYTNdraU2DseOJG5G0oQsyhQBFlczNyPA4Xxnyiu7wELkoa1v73+VcBuQX8NU9Mcmz3ifS
H0J+IlI5QNyrvDBzoLztqlSw47rJNgCKbD+cGZkyVguOnstXCE5YaDbSDuhuV9U+83tnXMQXcNqY
gcXFc7AqUEdOqfYr1Ou2McfhJET+cRRKQXLD/F5XU3je14NnQwIdmQMyiX4uenfCj3ZiK8cHLmjJ
PdNUDC7SbLncH4HqPZ7q9c38XUbd6FWOehsNRmIME6UvlCzGcwgeQlxq4xHSxGHyiaqrusKipmx9
2mom4MNXquNc/SrVkYWXt7vN8fs2x0Z8pjoqhSmDPE1wr0vjnMR1WYnsYN6v58/Mw9HNKPIVBH9Z
5oPp0WxRyDeqtFKa2VcweiXWhFhiI4bL/34WFq2UnbnQPIfW8ABjl3CRjtMhTpzMzhFhDawcQ13T
I9vTYzGQispHI42v9SaOtBUGgPnLATThVNXKsJ/VYo7g3xN4DHDSusehbkgzI1i2zS26nFw2frlh
NrN8YXe5vexgkJAutgiVYvHPjDTUWo+ByymiSBMgo4+TZWHlfeR1HsXZopuBIil5S0jNwq+V0Fob
Yu5xfm9Dw/PIi1crwQH/3ZG/2K4wTCj9zFXPf4yIulpQvn1PFe/SLiWIUwnwtzZCWugc7iabhGmY
LEKe9DUOY1G6TsMZUtWMr4bZ5lw9ns+15l3Kd9IQxx2l6OQX/sJd8npLR5sHfGhM973G7eSHQ+87
H6M0lhOzV2gA0h2UNClEh2Eewk0q4UBWU9FENE5M9szouXeyy/FhOKC3+WXhLyw6aN+meZ//5Aot
MR0VUy7LywR11gk6vNOLLuyi0pF3Kz2MwFKR3WX4j8meTHilevJ/KHlSDpJJNr6RFvMbocOJk0bx
P6lTLwySwxAUBkNEF2or4sTcIUIgVx0riacKzmc4Db2YY0DNbOr2AUuzVSJg7KHLOiKJc0fRlbTO
5NW4+4INgK2nEaa1HD2poVUqVA1GtSElSEne4w+D3RV++ESqHxphkJFVFrbEXcwm/Joka9oFOMuv
T8O8TH1hYKRsMU7xDPXlu7folpBt8wvLFeeM7Ur8z4imeTvzokIkRZ3vpiGOScr6fYhyzCfFTG/F
aI8tqlQNLMZnIiWMgIIIB7TVk382SVnhf2VmfSlM7lfNTYAiqrk0gof4U/C0HCgNIfyy2BZQccmw
meL3BEHw661PVHlrigwvypgTUNLGoGL9wobu8V0VuYLYmkNltmH4jcw1oFKcNT0SgeC/jotcLWhb
0W4/gAdjuKqEVcrkRvvdHHYpqvHOWM6THA6/pMwK6yeRIRkpNVLFuOjzifEQ7qfbwqFo2nNWyipm
0DU+N3yfQNXbBtPaFbGPPStOcNN8nkflHgL+AXIfAur+jkSNlqDTEqZLyfCy4wT+I3JKq6prvrW7
JdsQGixIhZ2nhFJoGTlohe6m51rVSTWy9ORt7IJkwexGhTSzylQyaify/rMO/4Pcs89nKDYT1PPS
dL9+ryGY7JU8g4bmMVMhq63lr9YOgTdm/wVbWuz1G+ornZLHCKpZxUQqWPCbFpuU0XJG0AuxwYyc
Dqbwg7iiNQcAcR52v3KUKSBLT7DdyMsrKb1LFzteBYUl2rjb2VoDhxg99Jn921xgPZnjnJfjPK+/
SQotsJJleCkxsLODAQEnWebGOlMyPBDf3W6MhvSFw+lyS+U32KX2MxmcDrJ8v7/Y6g4sgQijFS8D
Sl31q6MoluwxjwbDecEhn0awpp19hOfJiZ456flEq2a4OsXO/PA8i5D++La5HaxSgEAK+sseeS0C
kp8yoiZb80A/5c87L9ycc9JQLhx2qYxuxfkdwXB5oEcqw7+noDS9X5UHLzv32cG1LHTmnwu5kB6F
0w6rm0bMaKQt9PXuJlwxgCR7atr4WiutHtvWEHtVqI9vvHhZfqeslgPuWJrRn38ZpK8/8tUGfAWp
XP6JxDWmMSkwpVSucootUfr5IONtcf7sEIyZ+pQnbkOhWYtOXyjLij/S4qIOBVySdZeZzOjV0gJb
7DmoxHNjpE6k3cZBNvn3PHPkHI8YqLfYlbIzsgauXbb55SLKOoRdkn6rumQq/fYFyV6WUFZDAE8Q
7rwQjHIikirB0U+C3d3ZaZlbAXA517qV/Ey/yonxLH4tDkkfCba1e2KV5RTy+H7P+L8u2mfDUWq3
AEXGfIV0+A5MAicg79I+7edH/fdvH67UNTETRe25NcZ5WxThKHjPmudV0j4TafxxfV+iv0wp6Zzz
aI9WFNm3AtVGCNNgM8drDmUh+UGBpyuiQZMGOhBoe0xXUvUXFn7EvI9a3SDtpiwyxziDvVBxmHBH
6IzE9yMPI7j1T6J+V3vOwb2Fq9zBsDLgCEO4UurH521k0FwYD33XdsDTtvWcVsUKdfs+iCqnOf4o
dE1aJzpZWzeOeuogYs0kf1foaI7HUjV5VNCAEKxPwaDum75+lDlYBwbF1A0sG4SakWbgWLnu8pQE
D+uWZL3EyTcDIqC8fCgldG7gAlyQtkt5kaeUTpZBiVGf9RZu5abXu2nNFDdm/txvuSJc9b5YeKah
sJp5mQrT8iP49HNAKUvifmHkckjIhTnkUrH81UDa23SH3mAGtjXRkiw4UpT66Ucl8eoTiK0zTY4i
/SZi5r95bhfpaybSUeNVYQbpm7B9RmE1U4ws3mCq6WGVpG8/ZyvQ3llWyw3tRspAtSED0FYcUNZt
Pik0RiULLvReFC+GuzcVqLR6upIQ0EbUylLl5Xj8j89VZaj3S4tO923hDDagBR0rAgb3DPwM/YIe
JTLDR385L8bPhxFWT9YBoH3bTwoViF6qB2I1U+aAm6Um1lJIeZM3pD0TKG1Ab7oRiXYcny7wTdvZ
aNM3mpOtNIGeuTDpVx6E5vcPyfz8Dr2Bzf6QcF6E7mwCjKBpziDB7SjDUJjdhDov7YY1HedTQXQi
KcQ+AANi8epe5AzfsSTyV0Ip1sGKEk+PT7kslNAckaGKsrCM2bMIEUP5MTidxVTsAgvSwKgZX92k
57NDos9n+RmqFzuvt04VdYnzdhYZ88J7FpsLJSpTa9W1xbQ/muWXj0kg+bpCXJIw4EtlWJOKdkEG
nAU/J/BiVtF3AQtext1YsTDaN12XT4rp8jw4afmT5ki51lzzy1I3pXE6OjlpwGhbsgC6wSwMzwXA
COukxmjlM7quqDYZPG0WkgYfjf0o8FNwC9hLbiO5PA9/k58vyON0gB0uZ618Knms0H6hpC+KLxMr
togdOrNshBNIO6sshFm7vpOILsofqpInROw5/mfmOFrtxCyOw2puW118phnGp5DzcEkqSCdMQsjj
NchStSCul4nI/XdxstO+sE4eOvqaM3Hva5zRjkpr/oZ9IBe0qP7JssXqRHw0nZHvPEr1cON3GsfN
g58pqgjfkrWCyLXKkJK5bTTDRRolD8P7fSpIubOiqDjcK9Dlhs2YKoA/pYgmbPXcV87jE2LouLJT
O7Rqlmnj5K28xrQOThxkOuxzZX9SW0FVx7+LQZqBK37yBtgaZSCh+tbHyvhD9Y7X+mPBNDpXXXEf
0KSQkucFpsntlsEBTdBBEOvFztQIOWrM+8y1Qm5w9VZlhWt1Hc1ms/meTRCX+IDZsyZl8GMWcO3i
hU7aJttQDr3vyWAJiDJFjJWpd2GEjaupzEiKmXnrhgscHJ7U8aU9mtWGU17U8DT3MB+qQ6sSJQkR
O8iy/jckbOkFkZDEPIBgoWnYunzESXHhGbTbI6FfOtrnBYMjMM81Lz3QwSlV0HXEbmbRaC1Rrd6q
dBqhzhbk6aNZ6KTaQFK3ZQsqKYx0i7DP9eay5Rj0sJR8gEq4bEs2Up+b1nTscFRjPLjn1IZbBsof
tXT9dy/+E0qwqg+5ufBFT2KQYvgEapmM9TO5D5kGmkeky1zInlDnm8VVKq6HnAw2+4RRm9fQYmTh
Etm2oIPQbTk6aeJ9uDPlq3/mIjRhPu4eRiOThhxxK21flrurQS2yZMFvIz6ZRZHoeb/NeDjZAsbA
z9wOWvgo+uRgiLdt5DJ1V0h71rBuREDzLov3XMnmmwtiSO+xr5oQ4rfi2d7nqbwVdYXunIESVuae
ncmFRw92Vh87p9YYbyr9ga8mZ0DR1wYOGrdHKrfmVEQpFsSUuh22s2oDrV8qzxa318N+PTS9bCZW
+Y6V5VOnoGPlqZ/y09Hbb/I9nSfbIvQKUmWtUdwMPrMU7PP188KoQ9Xpe09HfDBv7yQ+xuJrYAuG
ykgaEKaFzgrBdX1NOLSbWkk7xHNp0fdbn/YacPThOXitqBqpvwyGlWyWipjwQtpQV7GFrVS8sbML
sYdNr1/5g8Uf1A9SvnCtBk+RLiOAqYRY8xMvtIu/9eBYHgebRWiqg24GzSURDE5nciKEqVW27UJ9
Oj2FhZ5KS9jfojVs8/klV0M+M07n8v1ejZZV+RV7qoJjmNI5JLcqsGi/ZCwTUjtpnWStdBlmXmVC
pWkivVPr9owgzrPcqw7mXwlIHeqdYZypuOJsGU2RIw9djXiPC1IorOyx/Nu1lN44Bkrn+/1dHt9H
Da4cgH1HcpEBSN+o42P97hRGxpS2CiiCgrLipPUmC6D1wrd81W8Ds+RgEXe7TOkpK1b6LBEPKdFv
csI0cokSB1q7OPvB5wQ3JusKWka3qX3hIsymey4PxdY1lEWAf0Kzm0VWq7e2qwxYNc/Tu9Ixp+Bx
v4TUZ/UZ2HzvKQmOWTQxbEQ9rBi7J8tJUrTI/qPbeU1PtRP71SGDBLY6MnXUs5dZtXIPr0+9y/El
DjkAHP1OPIQSZ+9ubuVmBARDdm+Td3RSt24/dM0j/mSgVNuYhVxtBxJ3K3WgaJP+WLRTsAcRTzPH
BMIPS8zPgUodN/1PR7JCzCLU0v8nrrD3i9x7Fq6KdjGyKBLqbL89iUYIAh8uOJUDh2GjliWpCMs/
dbsnfcIFbydODqsF5lxCy5CPFKSdoe2xIh8uSCLtOx+9sTlq3G0V4pghTqN75TffkNT+7SqQSYpm
gldY79Q1ymjgbSdY+LoKJ624PuvwX7dWPSw9glrQi73prz/XAy8bnDi9HRD987Crj6agpx0JRNGE
sviuXr2Yr+tWOoR0mXnIwdGiBwUTdGOzYObtIWDQWxSkzu7X/DkgI0fABfVC0Zg6MgZdjGVBlJHv
plIhcuP8SxWNYPtx0DLr99XBgR+8Z5kqKKnP5F/etolk1TCb6tYRXVO7BFYkn7/2LasaVEI4/82K
QAnRUiczqINKreD43cytwJES44zBYqJanbvkWQg8sgThP3fho6gGQy4FMlY4A/3tuQw+HBr6XNBK
XNR4CBrTLzKTFdlYdhcMftG0EeXF/ya41U1J7yqFhSllo1Kow1O7D5TwG2MRDau7dc6+9F0Lt/ku
3wOZaoXLlm7oF4e2abga+x1+c34kkDttJ6v1oAGZ8ebQlPuBeMbJfPBT9QTOgYGa1pXusxKm6sf1
K/2q3CqNzgZwGFB7q1R2XvIIBgXPqCghI0ZwmDMqDvql5PMHqBrCY3fwztLUH3ILrikdOetvDG0n
EXKgw1uoPOJkICWkDTvULBs=
`protect end_protected
